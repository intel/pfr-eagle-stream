package gen_gpi_signals_pkg;

    localparam GPI_1_cc_RST_RSMRST_PLD_R_N_BIT_POS = 0;
    localparam GPI_1_cc_RST_SRST_BMC_PLD_R_N_BIT_POS = 1;
    localparam GPI_1_FM_ME_PFR_1_BIT_POS = 2;
    localparam GPI_1_FM_ME_PFR_2_BIT_POS = 3;
    localparam GPI_1_PLTRST_DETECTED_REARM_ACM_TIMER_BIT_POS = 4;
    localparam GPI_1_BMC_SPI_IBB_ACCESS_DETECTED_BIT_POS = 5;
    localparam GPI_1_FM_PFR_FORCE_RECOVERY_N_BIT_POS = 6;
    localparam GPI_1_HPFR_IN_BIT_POS = 7;
    localparam GPI_1_LEGACY_BIT_POS = 8;
    localparam GPI_1_HPFR_ACTIVE_BIT_POS = 9;
    localparam GPI_1_UNUSED_BITS_START_BIT_POS = 10;

endpackage
