/////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////
/*!

	\brief    <b>%Led Control  </b>
	\file     led_control.v
	\details    <b>This block is in charge of multiplexing the LED_CONTROL output </b>
                <b> various destinations as the STATUS LEDs, the 2 7-segment Displays </b>
                <b> the fan fault LEDs and the CPUs DIMM fault indications by using  </b>
                <b> separated select outputs for each destination </b>
                <b> We use the 2 dots (1 per display) to identify which post code we are posting </b>
                <b> 2 dots  --> MainFpga Postcodes </b>
                <b> 1 dot   --> PFR Postcodes </b>
                <b> no dots --> BIOS Postcodes </b>
                <b> Also, when the PLD_REV_N is asserted we display FPGA versions like this: </b>
                <b> 1 dot  --> MainFpga version </b>
                <b> 2 dots --> DebugFpga Postcodes </b>
								 
				
	\brief  <b> New block implementation</b> 
			$Date    : Sept 18, 2019 $
			$Author  : a.larios@intel.com $			
			Project  : Archer City RP
			Group    : BD
			   
	\copyright Intel Proprietary -- Copyright \htmlonly <script>document.write(new Date().getFullYear())</script> \endhtmlonly Intel -- All rights reserved */
////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////////



module led_control
  #(parameter MAINFPGAVER = 8'h01, DEBUGFPGAVER = 8'h01)
  (
    input       iClk,                             //%Clock input 
    input       iRst_n,                           //%Reset enable on Low

    input       iRstPltRst_n,                     //PLTRST_N signal comming from PCH (used to automatically switch from FPGA to BIOS postcodes in displays)

    input [7:0] iStatusLeds,                       //input to be reflected at status LEDs from BMC SGPIO when oStatusLedSel is asserted
    output reg  oStatusLedSel,                    //output generated by this module to select when STATUS LEDs should take into account the LED_CONTROL output pins

    input [7:0] iFpgaPostCode1,                   //Main Fpga postcode for 7-segment display 1 (MSB) before PLT_RST_N is deasserted (already encoded into 7-Seg Display)
    input [7:0] iFpgaPostCode2,                   //Main Fpga postcode for 7-segment display 2 (LSB) before PLT_RST_N is deasserted (already encoded into 7-seg Display)
    input [7:0] iBiosPostCode,                    //Port 80 post-codes from BIOS for the 2 7-Segment displays, after PLT_RST_N is deasserted
    input [7:0] iPFRPostCode,                    //PFR postcode to be displayed on 7-segment display 1 (MSB), by asserting PFR override signal (overriding Fpga & BIOS post-codes)
    //input [6:0] iPFRPostCode2,                    //PFR postcode to be displayed on 7-segment display 2 (LSB), by asserting PFR override signal (overriding Fpga & BIOS post-codes)
    input       iPFROverride,                     //PRF override signal, if asserted, PRF postcode data is displayed in 7-segment displays, otherwise, FPGA or BIOS postcodes will be displayed depending on RST_PLTRST_N signal
    output reg  oPostCodeSel1_n,                  //to latch LED_CONTROL outputs into the 7-segment display1 (MSB) (active low)
    output reg  oPostCodeSel2_n,                  //to latch LED_CONTROL outputs into the 7-segment display2 (LSB) (active low)

    input [7:0] iLedFanFault,                     //input to be reflected at FAN FAULT LEDs, latched into LED_CONTROL when oLedFanFaultSel is asserted
    output reg  oLedFanFaultSel_n,                //output to latch LED_CONTROL outputs into Fan Fault LEDs (active low)

    input [7:0] iLedCpu0DimmCh1Fault,               //input for the Cpu0 Dimms 1&2 CH 1-4 Fault LEDs indications
    output reg  oLedCpu0DimmCh1FaultSel,            //to latch LED_CONTROL output into CPU0 Dimms 1&2 on CH 1-4 Fault LEDs
   
    input [7:0] iLedCpu0DimmCh5Fault,               //input for the Cpu0 Dimms 1&2 CH 5-8 Fault LEDs indications
    output reg  oLedCpu0DimmCh5FaultSel,            //to latch LED_CONTROL output into CPU0 Dimms 1&2 on CH 5-8 Fault LEDs
   
    input [7:0] iLedCpu1DimmCh1Fault,               //input for the Cpu1 Dimms 1&2 CH 1-4 Fault LEDs indications
    output reg  oLedCpu1DimmCh1FaultSel,            //to latch LED_CONTROL output into CPU1 Dimms 1&2 on CH 1-4 Fault LEDs
   
    input [7:0] iLedCpu1DimmCh5Fault,               //input for the Cpu1 Dimms 1&2 CH 5-8 Fault LEDs indications
    output reg  oLedCpu1DimmCh5FaultSel,            //to latch LED_CONTROL output into CPU1 Dimms 1&2 on CH 5-8 Fault LEDs
   

/* -----\/----- EXCLUDED -----\/-----
    input [6:0] iMainFpgaVer1,                    //Main Fpga Version (MSB) to be displayed in 7-segment display1 (MSB)
    input [6:0] iMainFpgaVer2,                    //Main Fpga Version (LSB) to be displayed in 7-segment display2 (MSB)4

    input [6:0] iDebugFpgaVer1,                   //Main Fpga Version (MSB) to be displayed in 7-segment display1 (MSB)
    input [6:0] iDebugFpgaVer2,                   //Main Fpga Version (LSB) to be displayed in 7-segment display2 (MSB)
 -----/\----- EXCLUDED -----/\----- */

    input       iPldRev_n,                        //when asserted (active low) will show Main/Debug FPGA versions in 7-Segment Displays 2&1
   
    output      [7:0] oLedControl                 //output of the mux to all LEDs resources
   );


   //////////////////////////////////
   //local params declarations
   ////////////////////////////////////////////////////////////////// 
   
   localparam INIT          = 4'd0;
   localparam DISPLAY1      = 4'd1;
   localparam DISPLAY1_D    = 4'd2;
   localparam DISPLAY2      = 4'd3;
   localparam DISPLAY2_D    = 4'd4;
   localparam STATUSLEDS    = 4'd5;
   localparam FANLEDS       = 4'd6;
   localparam CPU0DIMM1LEDS = 4'd7;
   localparam CPU0DIMM2LEDS = 4'd8;
   localparam CPU1DIMM1LEDS = 4'd9;
   localparam CPU1DIMM2LEDS = 4'd10;

   localparam ENDVERCNT = 9'd299;
   

   //////////////////////////////////
   //internal signals declarations
   ////////////////////////////////////////////////////////////////// 

   reg [3:0]  rLedFsm;              //FSM for the LED_CONTROL muxing
   reg [7:0]  rLedControl;          //to register LED_CONTROL before output
   reg        rVerFlag;             //when PLD_REV_N button is pressed, this signal will toggle evey 1 sec to switch from Main 2 Debug PLD versions
   reg [8:0]  rVerCnt;              //from the 3.33 msec clock we will cnt to get a 1 second delay to toggle rVerFlag, so we can mux the Main & Debug versions displayed while PLD_REV_N is asserted
   
   
   
   //////////////////////////////////
   //local function to decode from Hex to 7-Segment Display & LED
   ////////////////////////////////////////////////////////////////// 

   function [7:0] fDecoder;
      input  [6:0] iEncodedData;      //data to be decoded into BCD 7-segments for displays
      input        iDotSel;           //it indicates if we need to turn the displays dots or not (depending if it is data for MainFpga (0), BIOS (1), or PFR (2)
      
      begin
		 case (iEncodedData)            //Decoder from decimal to 7 Seg
		   7'd0:  fDecoder[6:0] = 7'b1000000; //0 -- 40h
		   7'd1:  fDecoder[6:0] = 7'b1111001; //1 -- 79h
		   7'd2:  fDecoder[6:0] = 7'b0100100; //2 -- 24h
		   7'd3:  fDecoder[6:0] = 7'b0110000; //3 -- 30h
		   7'd4:  fDecoder[6:0] = 7'b0011001; //4 -- 19h
		   7'd5:  fDecoder[6:0] = 7'b0010010; //5 -- 12h
		   7'd6:  fDecoder[6:0] = 7'b0000010; //6 -- 02h
		   7'd7:  fDecoder[6:0] = 7'b1111000; //7 -- 78h
		   7'd8:  fDecoder[6:0] = 7'b0000000; //8 -- 00h
		   7'd9:  fDecoder[6:0] = 7'b0010000; //9 -- 10h
		   7'd10: fDecoder[6:0] = 7'b0001000; //A -- 08h
		   7'd11: fDecoder[6:0] = 7'b0000011; //b -- 03h
		   7'd12: fDecoder[6:0] = 7'b1000110; //C -- 46h
		   7'd13: fDecoder[6:0] = 7'b0100001; //d -- 21h
		   7'd14: fDecoder[6:0] = 7'b0000110; //E -- 06h
		   7'd15: fDecoder[6:0] = 7'b0001110; //F -- 0Eh
		   7'd16: fDecoder[6:0] = 7'b0111111; //- -- 3Fh
		   default: 
			 fDecoder[6:0] = 7'b1111111; //ALL OFF
         endcase // case (encoded_data)

         fDecoder[7] = iDotSel;
      end
   endfunction // decoder
   

   //////////////////////////////////
   //FSM for the LED_CONTROL muxing 
   ////////////////////////////////////////////////////////////////// 

   always @(posedge iClk)
     begin
        if (~iRst_n)
          begin
             rLedFsm <= INIT;
             oStatusLedSel <= 1'b0;    //active high
             
             oPostCodeSel1_n <= 1'b1;  //active low
             oPostCodeSel2_n <= 1'b1;  //active low
             
             oLedFanFaultSel_n <= 1'b1;  //active low
             
             oLedCpu0DimmCh1FaultSel <= 1'b0;  //active high
             oLedCpu0DimmCh5FaultSel <= 1'b0;  //active high
             oLedCpu1DimmCh1FaultSel <= 1'b0;  //active high
             oLedCpu1DimmCh5FaultSel <= 1'b0;  //active high

             rVerFlag <= 1'b0;
             rVerCnt <= 9'h0;
             
          end // if (~iRst_n)
        else
          begin

             //this will generate a 1-sec toggling signal to swith from main to debug fpga versions in the display when the PLD_REV_N is asserted
             if (~iPldRev_n)
               begin
                  if (rVerCnt == ENDVERCNT)
                    begin
                       rVerFlag <= ~rVerFlag;
                       rVerCnt <= 0;
                    end
                  else
                    rVerCnt <= rVerCnt + 1'b1;
               end
             else
               begin
                  rVerFlag <= 0;        //if PLD_REV_N is de-asserted, we go back to init state so always we start with the MainFPGA ver first, and then Debug, etc
                  rVerCnt <= 0;
               end

             case (rLedFsm)
               default: begin   //INIT && CPU1DIMM2LEDS
                  oLedCpu1DimmCh5FaultSel <= 1'b0;  //de-selecting CPU1 DIMM1 Fault LEDs
                  oPostCodeSel1_n <= 1'b0;      //enabling data to be in 7-Seg Display1 (MSB)

                  rLedFsm <= DISPLAY1;

                  if (~iPldRev_n)
                    begin
                       
                       if (rVerFlag == 1'b0)
                         rLedControl <= fDecoder({3'h0,MAINFPGAVER[7:4]},0);              //if PldRev_n button is pushed, it shows Main and Debg Fpga versions (middle dot ON)
                       else
                         rLedControl <= fDecoder({3'h0,DEBUGFPGAVER[7:4]},0);             //if PldRev_n button is pushed, it shows Main and Debg Fpga versions (middle dot ON)
                       
                    end
                  else
                    begin
                       if (iPFROverride == 1'b1)                                          //if PFROverride is asserted, select PFR postcodes over MainFPGA or BIOS
                         begin
                            rLedControl <= fDecoder({3'h0,iPFRPostCode[7:4]},1);          //middle dot OFF
                         end
                       else
                         begin
                            if (iRstPltRst_n == 1'b0)                                     //if not PFROverride and PLT RST is yet asserted, do MainFPGA postcodes
                              begin
                                 rLedControl <= iFpgaPostCode1;                           //middle dot ON
                              end
                            else
                              begin                                                       //When PLT_RST is deasserted and no override asserted, do BIOS post codes
                                 rLedControl <= fDecoder({3'h0,iBiosPostCode[7:4]},1);    //middle dot OFF
                              end
                         end // else: !if(iPFROverride == 1'b1)
                    end // else: !if(~iPldRev_n)
               end // case: default

               DISPLAY1:begin
                  rLedFsm <= DISPLAY1_D;                                                 //to give an extra cycle to Display1
               end
                 
               DISPLAY1_D: begin
                  rLedFsm <= DISPLAY2;
                  oPostCodeSel1_n <= 1'b1;      //disabling data for 7-Seg Display1 (MSB)
                  oPostCodeSel2_n <= 1'b0;      //enabling data to be in 7-Seg Display2 (LSB)

                  if (~iPldRev_n)
                    begin
                       
                       if (rVerFlag == 1'b0)
                         rLedControl <= fDecoder({3'h0,MAINFPGAVER[3:0]},1);              //if PldRev_n button is pushed, it shows Main and Debg Fpga versions (end dot OFF)
                       else
                         rLedControl <= fDecoder({3'h0,DEBUGFPGAVER[3:0]},0);             //if PldRev_n button is pushed, it shows Main and Debg Fpga versions (end dot ON)
                    end
                  else
                    begin
                       if (iPFROverride == 1'b1)                                          //if PFROverride is asserted, select PFR postcodes over MainFPGA or BIOS
                         begin
                            rLedControl <= fDecoder({3'h0,iPFRPostCode[3:0]},0);          //end dot ON
                         end
                       else
                         begin
                            if (iRstPltRst_n == 1'b0)                                     //if not PFROverride and PLT RST is yet asserted, do MainFPGA postcodes
                              begin
                                 rLedControl <= iFpgaPostCode2;                           //end dot ON
                              end
                            else
                              begin                                                       //When PLT_RST is deasserted and no override asserted, do BIOS post codes
                                 rLedControl <= fDecoder({3'h0,iBiosPostCode[3:0]},1);    //end dot OFF
                              end
                         end // else: !if(iPFROverride == 1'b1)
                    end // else: !if(~iPldRev_n)
               end // case: 7SEG1

               DISPLAY2:begin
                  rLedFsm <= DISPLAY2_D;                                                 //to give an extra cycle to Display2
               end

               DISPLAY2_D: begin
                  rLedFsm <= STATUSLEDS;
                  oPostCodeSel2_n <= 1'b1;       //de-selecting Display2 
                  oStatusLedSel <= 1'b1;         //selecting STATUS LEDs
                  
                  rLedControl <= iStatusLeds;    ////data coming from BMC SGPIO for Status LEDs
               end //case: 7SEG2

               STATUSLEDS: begin
                  oStatusLedSel <= 1'b0;         //de-selecting status LEDs
                  oLedFanFaultSel_n <= 1'b0;     //selecting fan-fault LEDs

                  rLedControl <= iLedFanFault;   //data coming from BMC SGPIO for fan fault indications

                  rLedFsm <= FANLEDS;            
               end //case: STATUSLEDS

               FANLEDS: begin
                  oLedFanFaultSel_n <= 1'b1;      //de-selecting fan-fault LEDs
                  oLedCpu0DimmCh1FaultSel <= 1'b1;  //selecting CPU0 DIMM1 Fault LEDs
                  
                 
                  rLedControl <= iLedCpu0DimmCh1Fault;   //data coming from BMC SGPIO for CPU0 DIMM1 Fault indications 
               
                  rLedFsm <= CPU0DIMM1LEDS;
               end //case: FANLEDS

               CPU0DIMM1LEDS: begin
                  oLedCpu0DimmCh1FaultSel <= 1'b0;  //de-selecting CPU0 DIMM1 Fault LEDs
                  oLedCpu0DimmCh5FaultSel <= 1'b1;  //selecting CPU0 DIMM2 Fault LEDs
                  
                 
                  rLedControl <= iLedCpu0DimmCh5Fault;   //data coming from BMC SGPIO for CPU0 DIMM2 Fault indications 
               
                  rLedFsm <= CPU0DIMM2LEDS;
               end //case: CPU0DIMM1LEDS

               CPU0DIMM2LEDS: begin
                  oLedCpu0DimmCh5FaultSel <= 1'b0;  //de-selecting CPU0 DIMM2 Fault LEDs
                  oLedCpu1DimmCh1FaultSel <= 1'b1;  //selecting CPU1 DIMM1 Fault LEDs
                  
                 
                  rLedControl <= iLedCpu1DimmCh1Fault;   //data coming from BMC SGPIO for CPU0 DIMM2 Fault indications 
               
                  rLedFsm <= CPU1DIMM1LEDS;
               end //case: CPU0DIMM2LEDS

               CPU1DIMM1LEDS: begin
                  oLedCpu1DimmCh1FaultSel <= 1'b0;  //de-selecting CPU1 DIMM1 Fault LEDs
                  oLedCpu1DimmCh5FaultSel <= 1'b1;  //selecting CPU1 DIMM2 Fault LEDs
                  
                 
                  rLedControl <= iLedCpu1DimmCh5Fault;   //data coming from BMC SGPIO for CPU0 DIMM2 Fault indications 
               
                  rLedFsm <= CPU1DIMM2LEDS;
               end //case: CPU1DIMM1LEDS
          
             endcase // case (rLedFsm)
             
                  
          end // else: !if(~iRst_n)
        

     end // always @ (posedge iClk)
   
   //////////////////////////////////
   //output assingments
   ////////////////////////////////////////////////////////////////// 

   assign oLedControl = rLedControl;
   

endmodule // led_control
