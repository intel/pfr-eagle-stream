wire FAN_BMC_PWM_R;
wire FM_ME_AUTHN_FAIL;
wire FM_ME_BT_DONE;
wire FM_PFR_DSW_PWROK_N;
wire FM_PFR_FORCE_RECOVERY_N;
wire FM_PFR_ON_R;
wire FM_PFR_POSTCODE_SEL_N;
wire FM_PFR_RNDGEN_AUX;
wire FM_PFR_SLP_SUS_EN_R_N;
wire FM_PFR_TM1_HOLD_N;
wire FM_SPI_PFR_BMC_BT_MASTER_SEL_R;
wire FM_SPI_PFR_PCH_MASTER_SEL_R;
wire FP_ID_LED_N;
wire FP_ID_LED_PFR_N;
wire FP_LED_STATUS_AMBER_N;
wire FP_LED_STATUS_AMBER_PFR_N;
wire FP_LED_STATUS_GREEN_N;
wire FP_LED_STATUS_GREEN_PFR_N;
wire LED_CONTROL_0;
wire LED_CONTROL_1;
wire LED_CONTROL_2;
wire LED_CONTROL_3;
wire LED_CONTROL_4;
wire LED_CONTROL_5;
wire LED_CONTROL_6;
wire LED_CONTROL_7;
wire RST_PFR_EXTRST_R_N;
wire RST_PFR_OVR_RTC_R;
wire RST_PFR_OVR_SRTC_R;
wire RST_PLTRST_PLD_N;
wire RST_SPI_PFR_BMC_BOOT_N;
wire RST_SPI_PFR_PCH_N;
wire SMB_BMC_HSBP_STBY_LVC3_SCL;
wire SMB_BMC_HSBP_STBY_LVC3_SDA;
wire SMB_PCH_PMBUS2_STBY_LVC3_SCL;
wire SMB_PCH_PMBUS2_STBY_LVC3_SDA;
wire SMB_PCIE_STBY_LVC3_B_SCL;
wire SMB_PCIE_STBY_LVC3_B_SDA;
wire SMB_PFR_HSBP_STBY_LVC3_SCL;
wire SMB_PFR_HSBP_STBY_LVC3_SDA;
wire SMB_PFR_PMB1_STBY_LVC3_SCL;
wire SMB_PFR_PMB1_STBY_LVC3_SDA;
wire SMB_PFR_PMBUS2_STBY_LVC3_R_SCL;
wire SMB_PFR_PMBUS2_STBY_LVC3_R_SDA;
wire SMB_PFR_RFID_STBY_LVC3_SCL;
wire SMB_PFR_RFID_STBY_LVC3_SDA;
wire SMB_PMBUS_SML1_STBY_LVC3_SCL;
wire SMB_PMBUS_SML1_STBY_LVC3_SDA;
wire SMB_S3M_CPU0_SCL_LVC1;
wire SMB_S3M_CPU0_SDA_LVC1;
wire SPI_BMC_BOOT_CS_N;
wire SPI_BMC_BT_MUXED_MON_CLK;
wire SPI_BMC_BT_MUXED_MON_IO2;
wire SPI_BMC_BT_MUXED_MON_IO3;
wire SPI_BMC_BT_MUXED_MON_MISO;
wire SPI_BMC_BT_MUXED_MON_MOSI;
wire SPI_PCH_CS1_N;
wire SPI_PCH_MUXED_MON_CLK;
wire SPI_PCH_MUXED_MON_IO0;
wire SPI_PCH_MUXED_MON_IO1;
wire SPI_PCH_MUXED_MON_IO2;
wire SPI_PCH_MUXED_MON_IO3;
wire SPI_PCH_PFR_CS0_N;
wire SPI_PCH_TPM_CS_N;
wire SPI_PFR_BMC_BOOT_R_IO2;
wire SPI_PFR_BMC_BOOT_R_IO3;
wire SPI_PFR_BMC_BT_SECURE_CS_R_N;
wire SPI_PFR_BMC_FLASH1_BT_CLK;
wire SPI_PFR_BMC_FLASH1_BT_MISO;
wire SPI_PFR_BMC_FLASH1_BT_MOSI;
wire SPI_PFR_PCH_R_CLK;
wire SPI_PFR_PCH_R_IO0;
wire SPI_PFR_PCH_R_IO1;
wire SPI_PFR_PCH_R_IO2;
wire SPI_PFR_PCH_R_IO3;
wire SPI_PFR_PCH_SECURE_CS0_R_N;
wire SPI_PFR_PCH_SECURE_CS1_N;
wire SPI_PFR_TPM_CS_R2_N;
wire RST_RSMRST_PLD_R_N;
wire RST_SRST_BMC_PLD_R_N;
wire FM_POSTLED_SEL;
wire FM_POST_7SEG1_SEL_N;
wire FM_POST_7SEG2_SEL_N;



top dut
(
    .CLK_25M_OSC_MAIN_FPGA(CLK_25M_OSC_MAIN_FPGA),
    .FAN_BMC_PWM_R(FAN_BMC_PWM_R),
    .FM_AUX_SW_EN(common_core_if_bfm.FM_AUX_SW_EN),
    .FM_BMC_NMI_PCH_EN(common_core_if_bfm.FM_BMC_NMI_PCH_EN),
    .FM_BMC_ONCTL_N_PLD(common_core_if_bfm.FM_BMC_ONCTL_N_PLD),
    .FM_BMC_PFR_PWRBTN_OUT_R_N(common_core_if_bfm.FM_BMC_PFR_PWRBTN_OUT_R_N),
    .FM_BMC_PWRBTN_OUT_N(common_core_if_bfm.FM_BMC_PWRBTN_OUT_N),
    .FM_CPU0_INTR_PRSNT(common_core_if_bfm.FM_CPU0_INTR_PRSNT),
    .FM_CPU0_PKGID0(common_core_if_bfm.FM_CPU0_PKGID0),
    .FM_CPU0_PKGID1(common_core_if_bfm.FM_CPU0_PKGID1),
    .FM_CPU0_PKGID2(common_core_if_bfm.FM_CPU0_PKGID2),
    .FM_CPU0_PROC_ID0(common_core_if_bfm.FM_CPU0_PROC_ID0),
    .FM_CPU0_PROC_ID1(common_core_if_bfm.FM_CPU0_PROC_ID1),
    .FM_CPU0_SKTOCC_LVT3_PLD_N(common_core_if_bfm.FM_CPU0_SKTOCC_LVT3_PLD_N),
    .FM_CPU1_PKGID0(common_core_if_bfm.FM_CPU1_PKGID0),
    .FM_CPU1_PKGID1(common_core_if_bfm.FM_CPU1_PKGID1),
    .FM_CPU1_PKGID2(common_core_if_bfm.FM_CPU1_PKGID2),
    .FM_CPU1_PROC_ID0(common_core_if_bfm.FM_CPU1_PROC_ID0),
    .FM_CPU1_PROC_ID1(common_core_if_bfm.FM_CPU1_PROC_ID1),
    .FM_CPU1_SKTOCC_LVT3_PLD_N(common_core_if_bfm.FM_CPU1_SKTOCC_LVT3_PLD_N),
    .FM_DIMM_12V_CPS_S5_N(common_core_if_bfm.FM_DIMM_12V_CPS_S5_N),
    .FM_FORCE_PWRON_LVC3(common_core_if_bfm.FM_FORCE_PWRON_LVC3),
    .FM_ME_AUTHN_FAIL(FM_ME_AUTHN_FAIL),
    .FM_ME_BT_DONE(FM_ME_BT_DONE),
    .FM_P1V0_BMC_AUX_EN(common_core_if_bfm.FM_P1V0_BMC_AUX_EN),
    .FM_P1V05_PCH_AUX_EN(common_core_if_bfm.FM_P1V05_PCH_AUX_EN),
    .FM_P1V2_BMC_AUX_EN(common_core_if_bfm.FM_P1V2_BMC_AUX_EN),
    .FM_P2V5_BMC_AUX_EN(common_core_if_bfm.FM_P2V5_BMC_AUX_EN),
    .FM_P5V_EN(common_core_if_bfm.FM_P5V_EN),
    .FM_PCH_P1V8_AUX_EN(common_core_if_bfm.FM_PCH_P1V8_AUX_EN),
    .FM_PCH_PRSNT_N(common_core_if_bfm.FM_PCH_PRSNT_N),
    .FM_PFR_DSW_PWROK_N(FM_PFR_DSW_PWROK_N),
    .FM_PFR_FORCE_RECOVERY_N(FM_PFR_FORCE_RECOVERY_N),
    .FM_PFR_MUX_OE_CTL_PLD(common_core_if_bfm.FM_PFR_MUX_OE_CTL_PLD),
    .FM_PFR_ON_R(FM_PFR_ON_R),
    .FM_PFR_POSTCODE_SEL_N(FM_PFR_POSTCODE_SEL_N),
    .FM_PFR_RNDGEN_AUX(FM_PFR_RNDGEN_AUX),
    .FM_PFR_SLP_SUS_EN_R_N(FM_PFR_SLP_SUS_EN_R_N),
    .FM_PFR_TM1_HOLD_N(FM_PFR_TM1_HOLD_N),
    .FM_PLD_CLK_25M_R_EN(common_core_if_bfm.FM_PLD_CLK_25M_R_EN),
    .FM_PLD_CLKS_DEV_R_EN(common_core_if_bfm.FM_PLD_CLKS_DEV_R_EN),
    .FM_PLD_HEARTBEAT_LVC3(common_core_if_bfm.FM_PLD_HEARTBEAT_LVC3),
    .FM_PLD_REV_N(common_core_if_bfm.FM_PLD_REV_N),
    .FM_PS_EN_PLD_R(common_core_if_bfm.FM_PS_EN_PLD_R),
    .FM_PVCCD_HV_CPU0_EN(common_core_if_bfm.FM_PVCCD_HV_CPU0_EN),
    .FM_PVCCD_HV_CPU1_EN(common_core_if_bfm.FM_PVCCD_HV_CPU1_EN),
    .FM_PVCCFA_EHV_CPU0_R_EN(common_core_if_bfm.FM_PVCCFA_EHV_CPU0_R_EN),
    .FM_PVCCFA_EHV_CPU1_R_EN(common_core_if_bfm.FM_PVCCFA_EHV_CPU1_R_EN),
    .FM_PVCCFA_EHV_FIVRA_CPU0_R_EN(common_core_if_bfm.FM_PVCCFA_EHV_FIVRA_CPU0_R_EN),
    .FM_PVCCFA_EHV_FIVRA_CPU1_R_EN(common_core_if_bfm.FM_PVCCFA_EHV_FIVRA_CPU1_R_EN),
    .FM_PVCCIN_CPU0_R_EN(common_core_if_bfm.FM_PVCCIN_CPU0_R_EN),
    .FM_PVCCIN_CPU1_R_EN(common_core_if_bfm.FM_PVCCIN_CPU1_R_EN),
    .FM_PVCCINFAON_CPU0_R_EN(common_core_if_bfm.FM_PVCCINFAON_CPU0_R_EN),
    .FM_PVCCINFAON_CPU1_R_EN(common_core_if_bfm.FM_PVCCINFAON_CPU1_R_EN),
    .FM_PVNN_MAIN_CPU0_EN(common_core_if_bfm.FM_PVNN_MAIN_CPU0_EN),
    .FM_PVNN_MAIN_CPU1_EN(common_core_if_bfm.FM_PVNN_MAIN_CPU1_EN),
    .FM_PVNN_PCH_AUX_EN(common_core_if_bfm.FM_PVNN_PCH_AUX_EN),
    .FM_PVPP_HBM_CPU0_EN(common_core_if_bfm.FM_PVPP_HBM_CPU0_EN),
    .FM_PVPP_HBM_CPU1_EN(common_core_if_bfm.FM_PVPP_HBM_CPU1_EN),
    .FM_RST_PERST_BIT0(common_core_if_bfm.FM_RST_PERST_BIT0),
    .FM_RST_PERST_BIT1(common_core_if_bfm.FM_RST_PERST_BIT1),
    .FM_RST_PERST_BIT2(common_core_if_bfm.FM_RST_PERST_BIT2),
    .FM_SLP_SUS_RSM_RST_N(common_core_if_bfm.FM_SLP_SUS_RSM_RST_N),
    .FM_SLPS3_PLD_N(common_core_if_bfm.FM_SLPS3_PLD_N),
    .FM_SLPS4_PLD_N(common_core_if_bfm.FM_SLPS4_PLD_N),
    .FM_SPI_PFR_BMC_BT_MASTER_SEL_R(FM_SPI_PFR_BMC_BT_MASTER_SEL_R),
    .FM_SPI_PFR_PCH_MASTER_SEL_R(FM_SPI_PFR_PCH_MASTER_SEL_R),
    .FM_SX_SW_P12V_R_EN(common_core_if_bfm.FM_SX_SW_P12V_R_EN),
    .FM_SX_SW_P12V_STBY_R_EN(common_core_if_bfm.FM_SX_SW_P12V_STBY_R_EN),
    .FM_SYS_THROTTLE_R_N(common_core_if_bfm.FM_SYS_THROTTLE_R_N),
    .FM_THERMTRIP_DLY_LVC1_R_N(common_core_if_bfm.FM_THERMTRIP_DLY_LVC1_R_N),
    .FP_ID_LED_N(FP_ID_LED_N),
    .FP_ID_LED_PFR_N(FP_ID_LED_PFR_N),
    .FP_LED_STATUS_AMBER_N(FP_LED_STATUS_AMBER_N),
    .FP_LED_STATUS_AMBER_PFR_N(FP_LED_STATUS_AMBER_PFR_N),
    .FP_LED_STATUS_GREEN_N(FP_LED_STATUS_GREEN_N),
    .FP_LED_STATUS_GREEN_PFR_N(FP_LED_STATUS_GREEN_PFR_N),
    .H_CPU0_MEMHOT_IN_LVC1_R_N(common_core_if_bfm.H_CPU0_MEMHOT_IN_LVC1_R_N),
    .H_CPU0_MEMHOT_OUT_LVC1_N(common_core_if_bfm.H_CPU0_MEMHOT_OUT_LVC1_N),
    .H_CPU0_MEMTRIP_LVC1_N(common_core_if_bfm.H_CPU0_MEMTRIP_LVC1_N),
    .H_CPU0_MON_FAIL_PLD_LVC1_N(common_core_if_bfm.H_CPU0_MON_FAIL_PLD_LVC1_N),
    .H_CPU0_PROCHOT_LVC1_R_N(common_core_if_bfm.H_CPU0_PROCHOT_LVC1_R_N),
    .H_CPU0_THERMTRIP_LVC1_N(common_core_if_bfm.H_CPU0_THERMTRIP_LVC1_N),
    .H_CPU1_MEMHOT_IN_LVC1_R_N(common_core_if_bfm.H_CPU1_MEMHOT_IN_LVC1_R_N),
    .H_CPU1_MEMHOT_OUT_LVC1_N(common_core_if_bfm.H_CPU1_MEMHOT_OUT_LVC1_N),
    .H_CPU1_MEMTRIP_LVC1_N(common_core_if_bfm.H_CPU1_MEMTRIP_LVC1_N),
    .H_CPU1_MON_FAIL_PLD_LVC1_N(common_core_if_bfm.H_CPU1_MON_FAIL_PLD_LVC1_N),
    .H_CPU1_PROCHOT_LVC1_R_N(common_core_if_bfm.H_CPU1_PROCHOT_LVC1_R_N),
    .H_CPU1_THERMTRIP_LVC1_N(common_core_if_bfm.H_CPU1_THERMTRIP_LVC1_N),
    .IRQ_CPU0_MEM_VRHOT_N(common_core_if_bfm.IRQ_CPU0_MEM_VRHOT_N),
    .IRQ_CPU0_VRHOT_N(common_core_if_bfm.IRQ_CPU0_VRHOT_N),
    .IRQ_CPU1_MEM_VRHOT_N(common_core_if_bfm.IRQ_CPU1_MEM_VRHOT_N),
    .IRQ_CPU1_VRHOT_N(common_core_if_bfm.IRQ_CPU1_VRHOT_N),
    .LED_CONTROL_0(LED_CONTROL_0),
    .LED_CONTROL_1(LED_CONTROL_1),
    .LED_CONTROL_2(LED_CONTROL_2),
    .LED_CONTROL_3(LED_CONTROL_3),
    .LED_CONTROL_4(LED_CONTROL_4),
    .LED_CONTROL_5(LED_CONTROL_5),
    .LED_CONTROL_6(LED_CONTROL_6),
    .LED_CONTROL_7(LED_CONTROL_7),
    .M_AB_CPU0_FPGA_RESET_R_N(common_core_if_bfm.M_AB_CPU0_FPGA_RESET_R_N),
    .M_AB_CPU0_RESET_N(common_core_if_bfm.M_AB_CPU0_RESET_N),
    .M_AB_CPU1_FPGA_RESET_R_N(common_core_if_bfm.M_AB_CPU1_FPGA_RESET_R_N),
    .M_AB_CPU1_RESET_N(common_core_if_bfm.M_AB_CPU1_RESET_N),
    .M_CD_CPU0_FPGA_RESET_R_N(common_core_if_bfm.M_CD_CPU0_FPGA_RESET_R_N),
    .M_CD_CPU0_RESET_N(common_core_if_bfm.M_CD_CPU0_RESET_N),
    .M_CD_CPU1_FPGA_RESET_R_N(common_core_if_bfm.M_CD_CPU1_FPGA_RESET_R_N),
    .M_CD_CPU1_RESET_N(common_core_if_bfm.M_CD_CPU1_RESET_N),
    .M_EF_CPU0_FPGA_RESET_R_N(common_core_if_bfm.M_EF_CPU0_FPGA_RESET_R_N),
    .M_EF_CPU0_RESET_N(common_core_if_bfm.M_EF_CPU0_RESET_N),
    .M_EF_CPU1_FPGA_RESET_R_N(common_core_if_bfm.M_EF_CPU1_FPGA_RESET_R_N),
    .M_EF_CPU1_RESET_N(common_core_if_bfm.M_EF_CPU1_RESET_N),
    .M_GH_CPU0_FPGA_RESET_R_N(common_core_if_bfm.M_GH_CPU0_FPGA_RESET_R_N),
    .M_GH_CPU0_RESET_N(common_core_if_bfm.M_GH_CPU0_RESET_N),
    .M_GH_CPU1_FPGA_RESET_R_N(common_core_if_bfm.M_GH_CPU1_FPGA_RESET_R_N),
    .M_GH_CPU1_RESET_N(common_core_if_bfm.M_GH_CPU1_RESET_N),
    .PWRGD_CPU0_LVC1_R(common_core_if_bfm.PWRGD_CPU0_LVC1_R),
    .PWRGD_CPU1_LVC1_R(common_core_if_bfm.PWRGD_CPU1_LVC1_R),
    .PWRGD_CPUPWRGD_LVC1(common_core_if_bfm.PWRGD_CPUPWRGD_LVC1),
    .PWRGD_DRAMPWRGD_CPU0_AB_R_LVC1(common_core_if_bfm.PWRGD_DRAMPWRGD_CPU0_AB_R_LVC1),
    .PWRGD_DRAMPWRGD_CPU0_CD_R_LVC1(common_core_if_bfm.PWRGD_DRAMPWRGD_CPU0_CD_R_LVC1),
    .PWRGD_DRAMPWRGD_CPU0_EF_R_LVC1(common_core_if_bfm.PWRGD_DRAMPWRGD_CPU0_EF_R_LVC1),
    .PWRGD_DRAMPWRGD_CPU0_GH_R_LVC1(common_core_if_bfm.PWRGD_DRAMPWRGD_CPU0_GH_R_LVC1),
    .PWRGD_DRAMPWRGD_CPU1_AB_R_LVC1(common_core_if_bfm.PWRGD_DRAMPWRGD_CPU1_AB_R_LVC1),
    .PWRGD_DRAMPWRGD_CPU1_CD_R_LVC1(common_core_if_bfm.PWRGD_DRAMPWRGD_CPU1_CD_R_LVC1),
    .PWRGD_DRAMPWRGD_CPU1_EF_R_LVC1(common_core_if_bfm.PWRGD_DRAMPWRGD_CPU1_EF_R_LVC1),
    .PWRGD_DRAMPWRGD_CPU1_GH_R_LVC1(common_core_if_bfm.PWRGD_DRAMPWRGD_CPU1_GH_R_LVC1),
    .PWRGD_FAIL_CPU0_AB_PLD(common_core_if_bfm.PWRGD_FAIL_CPU0_AB_PLD),
    .PWRGD_FAIL_CPU0_CD_PLD(common_core_if_bfm.PWRGD_FAIL_CPU0_CD_PLD),
    .PWRGD_FAIL_CPU0_EF_PLD(common_core_if_bfm.PWRGD_FAIL_CPU0_EF_PLD),
    .PWRGD_FAIL_CPU0_GH_PLD(common_core_if_bfm.PWRGD_FAIL_CPU0_GH_PLD),
    .PWRGD_FAIL_CPU1_AB_PLD(common_core_if_bfm.PWRGD_FAIL_CPU1_AB_PLD),
    .PWRGD_FAIL_CPU1_CD_PLD(common_core_if_bfm.PWRGD_FAIL_CPU1_CD_PLD),
    .PWRGD_FAIL_CPU1_EF_PLD(common_core_if_bfm.PWRGD_FAIL_CPU1_EF_PLD),
    .PWRGD_FAIL_CPU1_GH_PLD(common_core_if_bfm.PWRGD_FAIL_CPU1_GH_PLD),
    .PWRGD_P1V0_BMC_AUX(common_core_if_bfm.PWRGD_P1V0_BMC_AUX),
    .PWRGD_P1V05_PCH_AUX(common_core_if_bfm.PWRGD_P1V05_PCH_AUX),
    .PWRGD_P1V2_BMC_AUX(common_core_if_bfm.PWRGD_P1V2_BMC_AUX),
    .PWRGD_P1V2_MAX10_AUX_PLD_R(common_core_if_bfm.PWRGD_P1V2_MAX10_AUX_PLD_R),
    .PWRGD_P1V8_PCH_AUX_PLD(common_core_if_bfm.PWRGD_P1V8_PCH_AUX_PLD),
    .PWRGD_P2V5_BMC_AUX(common_core_if_bfm.PWRGD_P2V5_BMC_AUX),
    .PWRGD_P3V3(common_core_if_bfm.PWRGD_P3V3),
    .PWRGD_PCH_PWROK_R(common_core_if_bfm.PWRGD_PCH_PWROK_R),
    .PWRGD_PLT_AUX_CPU0_LVT3_R(common_core_if_bfm.PWRGD_PLT_AUX_CPU0_LVT3_R),
    .PWRGD_PLT_AUX_CPU1_LVT3_R(common_core_if_bfm.PWRGD_PLT_AUX_CPU1_LVT3_R),
    .PWRGD_PS_PWROK_PLD_R(common_core_if_bfm.PWRGD_PS_PWROK_PLD_R),
    .PWRGD_PVCCD_HV_CPU0(common_core_if_bfm.PWRGD_PVCCD_HV_CPU0),
    .PWRGD_PVCCD_HV_CPU1(common_core_if_bfm.PWRGD_PVCCD_HV_CPU1),
    .PWRGD_PVCCFA_EHV_CPU0(common_core_if_bfm.PWRGD_PVCCFA_EHV_CPU0),
    .PWRGD_PVCCFA_EHV_CPU1(common_core_if_bfm.PWRGD_PVCCFA_EHV_CPU1),
    .PWRGD_PVCCFA_EHV_FIVRA_CPU0(common_core_if_bfm.PWRGD_PVCCFA_EHV_FIVRA_CPU0),
    .PWRGD_PVCCFA_EHV_FIVRA_CPU1(common_core_if_bfm.PWRGD_PVCCFA_EHV_FIVRA_CPU1),
    .PWRGD_PVCCIN_CPU0(common_core_if_bfm.PWRGD_PVCCIN_CPU0),
    .PWRGD_PVCCIN_CPU1(common_core_if_bfm.PWRGD_PVCCIN_CPU1),
    .PWRGD_PVCCINFAON_CPU0(common_core_if_bfm.PWRGD_PVCCINFAON_CPU0),
    .PWRGD_PVCCINFAON_CPU1(common_core_if_bfm.PWRGD_PVCCINFAON_CPU1),
    .PWRGD_PVNN_MAIN_CPU0(common_core_if_bfm.PWRGD_PVNN_MAIN_CPU0),
    .PWRGD_PVNN_MAIN_CPU1(common_core_if_bfm.PWRGD_PVNN_MAIN_CPU1),
    .PWRGD_PVNN_PCH_AUX(common_core_if_bfm.PWRGD_PVNN_PCH_AUX),
    .PWRGD_PVPP_HBM_CPU0(common_core_if_bfm.PWRGD_PVPP_HBM_CPU0),
    .PWRGD_PVPP_HBM_CPU1(common_core_if_bfm.PWRGD_PVPP_HBM_CPU1),
    .PWRGD_SYS_PWROK_R(common_core_if_bfm.PWRGD_SYS_PWROK_R),
    .RST_CPU0_LVC1_R_N(common_core_if_bfm.RST_CPU0_LVC1_R_N),
    .RST_CPU1_LVC1_R_N(common_core_if_bfm.RST_CPU1_LVC1_R_N),
    .RST_DEDI_BUSY_PLD_N(common_core_if_bfm.RST_DEDI_BUSY_PLD_N),
    .RST_PLD_PCIE_CPU0_DEV_PERST_N(common_core_if_bfm.RST_PLD_PCIE_CPU0_DEV_PERST_N),
    .RST_PLD_PCIE_CPU1_DEV_PERST_N(common_core_if_bfm.RST_PLD_PCIE_CPU1_DEV_PERST_N),
    .RST_PLD_PCIE_PCH_DEV_PERST_N(common_core_if_bfm.RST_PLD_PCIE_PCH_DEV_PERST_N),
    .RST_PFR_EXTRST_R_N(RST_PFR_EXTRST_R_N),
    .RST_PFR_OVR_RTC_R(RST_PFR_OVR_RTC_R),
    .RST_PFR_OVR_SRTC_R(RST_PFR_OVR_SRTC_R),
    .RST_PLTRST_PLD_B_N(common_core_if_bfm.RST_PLTRST_PLD_B_N),
    .RST_PLTRST_PLD_N(RST_PLTRST_PLD_N),
    .RST_SPI_PFR_BMC_BOOT_N(RST_SPI_PFR_BMC_BOOT_N),
    .RST_SPI_PFR_PCH_N(RST_SPI_PFR_PCH_N),
    .SGPIO_BMC_CLK(common_core_if_bfm.SGPIO_BMC_CLK),
    .SGPIO_BMC_DIN_R(common_core_if_bfm.SGPIO_BMC_DIN_R),
    .SGPIO_BMC_DOUT(common_core_if_bfm.SGPIO_BMC_DOUT),
    .SGPIO_BMC_LD_N(common_core_if_bfm.SGPIO_BMC_LD_N),
    .SMB_BMC_HSBP_STBY_LVC3_SCL(SMB_BMC_HSBP_STBY_LVC3_SCL),
    .SMB_BMC_HSBP_STBY_LVC3_SDA(SMB_BMC_HSBP_STBY_LVC3_SDA),
    .SMB_PCH_PMBUS2_STBY_LVC3_SCL(SMB_PCH_PMBUS2_STBY_LVC3_SCL),
    .SMB_PCH_PMBUS2_STBY_LVC3_SDA(SMB_PCH_PMBUS2_STBY_LVC3_SDA),
    .SMB_PCIE_STBY_LVC3_B_SCL(SMB_PCIE_STBY_LVC3_B_SCL),
    .SMB_PCIE_STBY_LVC3_B_SDA(SMB_PCIE_STBY_LVC3_B_SDA),
    .SMB_PFR_HSBP_STBY_LVC3_SCL(SMB_PFR_HSBP_STBY_LVC3_SCL),
    .SMB_PFR_HSBP_STBY_LVC3_SDA(SMB_PFR_HSBP_STBY_LVC3_SDA),
    .SMB_PFR_PMB1_STBY_LVC3_SCL(SMB_PFR_PMB1_STBY_LVC3_SCL),
    .SMB_PFR_PMB1_STBY_LVC3_SDA(SMB_PFR_PMB1_STBY_LVC3_SDA),
    .SMB_PFR_PMBUS2_STBY_LVC3_R_SCL(SMB_PFR_PMBUS2_STBY_LVC3_R_SCL),
    .SMB_PFR_PMBUS2_STBY_LVC3_R_SDA(SMB_PFR_PMBUS2_STBY_LVC3_R_SDA),
    .SMB_PFR_RFID_STBY_LVC3_SCL(SMB_PFR_RFID_STBY_LVC3_SCL),
    .SMB_PFR_RFID_STBY_LVC3_SDA(SMB_PFR_RFID_STBY_LVC3_SDA),
    .SMB_PMBUS_SML1_STBY_LVC3_SCL(SMB_PMBUS_SML1_STBY_LVC3_SCL),
    .SMB_PMBUS_SML1_STBY_LVC3_SDA(SMB_PMBUS_SML1_STBY_LVC3_SDA),
    .SMB_S3M_CPU0_SCL_LVC1(common_core_if_bfm.SMB_S3M_CPU0_SCL_LVC1),
    .SMB_S3M_CPU0_SCL_LVC1(SMB_S3M_CPU0_SCL_LVC1),
    .SMB_S3M_CPU0_SDA_LVC1(common_core_if_bfm.SMB_S3M_CPU0_SDA_LVC1),
    .SMB_S3M_CPU0_SDA_LVC1(SMB_S3M_CPU0_SDA_LVC1),
    .SMB_S3M_CPU1_SCL_LVC1(common_core_if_bfm.SMB_S3M_CPU1_SCL_LVC1),
    .SMB_S3M_CPU1_SDA_LVC1(common_core_if_bfm.SMB_S3M_CPU1_SDA_LVC1),
    .SPI_BMC_BOOT_CS_N(SPI_BMC_BOOT_CS_N),
    .SPI_BMC_BT_MUXED_MON_CLK(SPI_BMC_BT_MUXED_MON_CLK),
    .SPI_BMC_BT_MUXED_MON_IO2(SPI_BMC_BT_MUXED_MON_IO2),
    .SPI_BMC_BT_MUXED_MON_IO3(SPI_BMC_BT_MUXED_MON_IO3),
    .SPI_BMC_BT_MUXED_MON_MISO(SPI_BMC_BT_MUXED_MON_MISO),
    .SPI_BMC_BT_MUXED_MON_MOSI(SPI_BMC_BT_MUXED_MON_MOSI),
    .SPI_PCH_CS1_N(SPI_PCH_CS1_N),
    .SPI_PCH_MUXED_MON_CLK(SPI_PCH_MUXED_MON_CLK),
    .SPI_PCH_MUXED_MON_IO0(SPI_PCH_MUXED_MON_IO0),
    .SPI_PCH_MUXED_MON_IO1(SPI_PCH_MUXED_MON_IO1),
    .SPI_PCH_MUXED_MON_IO2(SPI_PCH_MUXED_MON_IO2),
    .SPI_PCH_MUXED_MON_IO3(SPI_PCH_MUXED_MON_IO3),
    .SPI_PCH_PFR_CS0_N(SPI_PCH_PFR_CS0_N),
    .SPI_PCH_TPM_CS_N(SPI_PCH_TPM_CS_N),
    .SPI_PFR_BMC_BOOT_R_IO2(SPI_PFR_BMC_BOOT_R_IO2),
    .SPI_PFR_BMC_BOOT_R_IO3(SPI_PFR_BMC_BOOT_R_IO3),
    .SPI_PFR_BMC_BT_SECURE_CS_R_N(SPI_PFR_BMC_BT_SECURE_CS_R_N),
    .SPI_PFR_BMC_FLASH1_BT_CLK(SPI_PFR_BMC_FLASH1_BT_CLK),
    .SPI_PFR_BMC_FLASH1_BT_MISO(SPI_PFR_BMC_FLASH1_BT_MISO),
    .SPI_PFR_BMC_FLASH1_BT_MOSI(SPI_PFR_BMC_FLASH1_BT_MOSI),
    .SPI_PFR_PCH_R_CLK(SPI_PFR_PCH_R_CLK),
    .SPI_PFR_PCH_R_IO0(SPI_PFR_PCH_R_IO0),
    .SPI_PFR_PCH_R_IO1(SPI_PFR_PCH_R_IO1),
    .SPI_PFR_PCH_R_IO2(SPI_PFR_PCH_R_IO2),
    .SPI_PFR_PCH_R_IO3(SPI_PFR_PCH_R_IO3),
    .SPI_PFR_PCH_SECURE_CS0_R_N(SPI_PFR_PCH_SECURE_CS0_R_N),
    .SPI_PFR_PCH_SECURE_CS1_N(SPI_PFR_PCH_SECURE_CS1_N),
    .SPI_PFR_TPM_CS_R2_N(SPI_PFR_TPM_CS_R2_N),
    .RST_RSMRST_PLD_R_N(RST_RSMRST_PLD_R_N),
    .RST_SRST_BMC_PLD_R_N(RST_SRST_BMC_PLD_R_N),
    .FM_POSTLED_SEL(FM_POSTLED_SEL),
    .FM_CPU_CATERR_LVT3_R_N(common_core_if_bfm.FM_CPU_CATERR_LVT3_R_N),
    .FM_ADR_ACK_R(common_core_if_bfm.FM_ADR_ACK_R),
    .FM_ADR_COMPLETE(common_core_if_bfm.FM_ADR_COMPLETE),
    .FM_ADR_TRIGGER_N(common_core_if_bfm.FM_ADR_TRIGGER_N),
    .FM_BMC_CRASHLOG_TRIG_N(common_core_if_bfm.FM_BMC_CRASHLOG_TRIG_N),
    .FM_PCH_CRASHLOG_TRIG_R_N(common_core_if_bfm.FM_PCH_CRASHLOG_TRIG_R_N),
    .FM_PCH_PLD_GLB_RST_WARN_N(common_core_if_bfm.FM_PCH_PLD_GLB_RST_WARN_N),
    .FM_PMBUS_ALERT_B_EN(common_core_if_bfm.FM_PMBUS_ALERT_B_EN),
    .FM_THROTTLE_R_N(common_core_if_bfm.FM_THROTTLE_R_N),
    .H_CPU_CATERR_LVC1_R_N(common_core_if_bfm.H_CPU_CATERR_LVC1_R_N),
    .H_CPU_NMI_LVC1_R(common_core_if_bfm.H_CPU_NMI_LVC1_R),
    .IRQ_BMC_CPU_NMI(common_core_if_bfm.IRQ_BMC_CPU_NMI),
    .IRQ_PCH_CPU_NMI_EVENT_N(common_core_if_bfm.IRQ_PCH_CPU_NMI_EVENT_N),
    .IRQ_SML1_PMBUS_PLD_ALERT_N(common_core_if_bfm.IRQ_SML1_PMBUS_PLD_ALERT_N),
    .FM_CPU1_DIMM_CH1_4_FAULT_LED_SEL(common_core_if_bfm.FM_CPU1_DIMM_CH1_4_FAULT_LED_SEL),
    .FM_CPU1_DIMM_CH5_8_FAULT_LED_SEL(common_core_if_bfm.FM_CPU1_DIMM_CH5_8_FAULT_LED_SEL),
    .FM_CPU0_DIMM_CH1_4_FAULT_LED_SEL(common_core_if_bfm.FM_CPU0_DIMM_CH1_4_FAULT_LED_SEL),
    .FM_CPU0_DIMM_CH5_8_FAULT_LED_SEL(common_core_if_bfm.FM_CPU0_DIMM_CH5_8_FAULT_LED_SEL),
    .FM_POST_7SEG1_SEL_N(FM_POST_7SEG1_SEL_N),
    .FM_POST_7SEG2_SEL_N(FM_POST_7SEG2_SEL_N),
    .FM_FAN_FAULT_LED_SEL_R_N(common_core_if_bfm.FM_FAN_FAULT_LED_SEL_R_N),
    .H_CPU_ERR0_LVC1_R_N(common_core_if_bfm.H_CPU_ERR0_LVC1_R_N),
    .H_CPU_ERR1_LVC1_R_N(common_core_if_bfm.H_CPU_ERR1_LVC1_R_N),
    .H_CPU_ERR2_LVC1_R_N(common_core_if_bfm.H_CPU_ERR2_LVC1_R_N),
    .FM_CPU_ERR0_LVT3_N(common_core_if_bfm.FM_CPU_ERR0_LVT3_N),
    .FM_CPU_ERR1_LVT3_N(common_core_if_bfm.FM_CPU_ERR1_LVT3_N),
    .FM_CPU_ERR2_LVT3_N(common_core_if_bfm.FM_CPU_ERR2_LVT3_N),
    .FM_DIS_PS_PWROK_DLY(common_core_if_bfm.FM_DIS_PS_PWROK_DLY),
    .FM_HBM2_HBM3_VPP_SEL(common_core_if_bfm.FM_HBM2_HBM3_VPP_SEL),
    .PWRGD_S0_PWROK_CPU0_LVC1_R(common_core_if_bfm.PWRGD_S0_PWROK_CPU0_LVC1_R),
    .PWRGD_S0_PWROK_CPU1_LVC1_R(common_core_if_bfm.PWRGD_S0_PWROK_CPU1_LVC1_R),
    .SGPIO_DEBUG_PLD_CLK(common_core_if_bfm.SGPIO_DEBUG_PLD_CLK),
    .SGPIO_DEBUG_PLD_DOUT(common_core_if_bfm.SGPIO_DEBUG_PLD_DOUT),
    .SGPIO_DEBUG_PLD_LD(common_core_if_bfm.SGPIO_DEBUG_PLD_LD),
    .SGPIO_DEBUG_PLD_DIN(common_core_if_bfm.SGPIO_DEBUG_PLD_DIN),
    .FP_BMC_PWR_BTN_R2_N(common_core_if_bfm.FP_BMC_PWR_BTN_R2_N),
    .FM_VAL_BOARD_PRSNT_N(common_core_if_bfm.FM_VAL_BOARD_PRSNT_N),
    .FM_ADR_MODE0(common_core_if_bfm.FM_ADR_MODE0),
    .FM_ADR_MODE1(common_core_if_bfm.FM_ADR_MODE1),
    .IRQ_BMC_PCH_NMI(common_core_if_bfm.IRQ_BMC_PCH_NMI),
    .FM_S3M_CPU0_CPLD_CRC_ERROR(common_core_if_bfm.FM_S3M_CPU0_CPLD_CRC_ERROR),
    .FM_S3M_CPU1_CPLD_CRC_ERROR(common_core_if_bfm.FM_S3M_CPU1_CPLD_CRC_ERROR),
    .SGPIO_IDV_CLK_R(common_core_if_bfm.SGPIO_IDV_CLK_R),
    .SGPIO_IDV_DOUT_R(common_core_if_bfm.SGPIO_IDV_DOUT_R),
    .SGPIO_IDV_DIN_R(common_core_if_bfm.SGPIO_IDV_DIN_R),
    .SGPIO_IDV_LD_R_N(common_core_if_bfm.SGPIO_IDV_LD_R_N),
)



