
`timescale 1 ps / 1 ps
`default_nettype none

module recovery_top (
    input wire CLK_25M_OSC_MAIN_FPGA,
    output wire FAN_BMC_PWM_R,
    output wire FM_AUX_SW_EN,
    input wire FM_BMC_NMI_PCH_EN,
    input wire FM_BMC_ONCTL_N_PLD,
    output wire FM_BMC_PFR_PWRBTN_OUT_R_N,
    input wire FM_BMC_PWRBTN_OUT_N,
    input wire FM_CPU0_INTR_PRSNT,
    input wire FM_CPU0_PKGID0,
    input wire FM_CPU0_PKGID1,
    input wire FM_CPU0_PKGID2,
    input wire FM_CPU0_PROC_ID0,
    input wire FM_CPU0_PROC_ID1,
    input wire FM_CPU0_SKTOCC_LVT3_PLD_N,
    input wire FM_CPU1_PKGID0,
    input wire FM_CPU1_PKGID1,
    input wire FM_CPU1_PKGID2,
    input wire FM_CPU1_PROC_ID0,
    input wire FM_CPU1_PROC_ID1,
    input wire FM_CPU1_SKTOCC_LVT3_PLD_N,
    input wire FM_DIMM_12V_CPS_S5_N,
    input wire FM_FORCE_PWRON_LVC3,
    input wire FM_ME_AUTHN_FAIL,
    input wire FM_ME_BT_DONE,
    output wire FM_P1V0_BMC_AUX_EN,
    output wire FM_P1V05_PCH_AUX_EN,
    output wire FM_P1V2_BMC_AUX_EN,
    output wire FM_P2V5_BMC_AUX_EN,
    output wire FM_P5V_EN,
    output wire FM_PCH_P1V8_AUX_EN,
    input wire FM_PCH_PRSNT_N,
    output wire FM_PFR_DSW_PWROK_N,
    input wire FM_PFR_FORCE_RECOVERY_N,
    output wire FM_PFR_MUX_OE_CTL_PLD,
    output wire FM_PFR_ON_R,
    input wire FM_PFR_POSTCODE_SEL_N,
    output wire FM_PFR_RNDGEN_AUX,
    output wire FM_PFR_SLP_SUS_EN_R_N,
    input wire FM_PFR_TM1_HOLD_N,
    output wire FM_PLD_CLK_25M_R_EN,
    output wire FM_PLD_CLKS_DEV_R_EN,
    output wire FM_PLD_HEARTBEAT_LVC3,
    input wire FM_PLD_REV_N,
    output wire FM_PS_EN_PLD_R,
    output wire FM_PVCCD_HV_CPU0_EN,
    output wire FM_PVCCD_HV_CPU1_EN,
    output wire FM_PVCCFA_EHV_CPU0_R_EN,
    output wire FM_PVCCFA_EHV_CPU1_R_EN,
    output wire FM_PVCCFA_EHV_FIVRA_CPU0_R_EN,
    output wire FM_PVCCFA_EHV_FIVRA_CPU1_R_EN,
    output wire FM_PVCCIN_CPU0_R_EN,
    output wire FM_PVCCIN_CPU1_R_EN,
    output wire FM_PVCCINFAON_CPU0_R_EN,
    output wire FM_PVCCINFAON_CPU1_R_EN,
    output wire FM_PVNN_MAIN_CPU0_EN,
    output wire FM_PVNN_MAIN_CPU1_EN,
    output wire FM_PVNN_PCH_AUX_EN,
    output wire FM_PVPP_HBM_CPU0_EN,
    output wire FM_PVPP_HBM_CPU1_EN,
    input wire FM_RST_PERST_BIT0,
    input wire FM_RST_PERST_BIT1,
    input wire FM_RST_PERST_BIT2,
    input wire FM_SLP_SUS_RSM_RST_N,
    input wire FM_SLPS3_PLD_N,
    input wire FM_SLPS4_PLD_N,
    output wire FM_SPI_PFR_BMC_BT_MASTER_SEL_R,
    output wire FM_SPI_PFR_PCH_MASTER_SEL_R,
    output wire FM_SX_SW_P12V_R_EN,
    output wire FM_SX_SW_P12V_STBY_R_EN,
    output wire FM_SYS_THROTTLE_R_N,
    output wire FM_THERMTRIP_DLY_LVC1_R_N,
    input wire FP_ID_LED_N,
    output wire FP_ID_LED_PFR_N,
    input wire FP_LED_STATUS_AMBER_N,
    output wire FP_LED_STATUS_AMBER_PFR_N,
    input wire FP_LED_STATUS_GREEN_N,
    output wire FP_LED_STATUS_GREEN_PFR_N,
    output wire H_CPU0_MEMHOT_IN_LVC1_R_N,
    input wire H_CPU0_MEMHOT_OUT_LVC1_N,
    input wire H_CPU0_MEMTRIP_LVC1_N,
    input wire H_CPU0_MON_FAIL_PLD_LVC1_N,
    output wire H_CPU0_PROCHOT_LVC1_R_N,
    input wire H_CPU0_THERMTRIP_LVC1_N,
    output wire H_CPU1_MEMHOT_IN_LVC1_R_N,
    input wire H_CPU1_MEMHOT_OUT_LVC1_N,
    input wire H_CPU1_MEMTRIP_LVC1_N,
    input wire H_CPU1_MON_FAIL_PLD_LVC1_N,
    output wire H_CPU1_PROCHOT_LVC1_R_N,
    input wire H_CPU1_THERMTRIP_LVC1_N,
    input wire IRQ_CPU0_MEM_VRHOT_N,
    input wire IRQ_CPU0_VRHOT_N,
    input wire IRQ_CPU1_MEM_VRHOT_N,
    input wire IRQ_CPU1_VRHOT_N,
    output wire LED_CONTROL_0,
    output wire LED_CONTROL_1,
    output wire LED_CONTROL_2,
    output wire LED_CONTROL_3,
    output wire LED_CONTROL_4,
    output wire LED_CONTROL_5,
    output wire LED_CONTROL_6,
    output wire LED_CONTROL_7,
    output wire M_AB_CPU0_FPGA_RESET_R_N,
    input wire M_AB_CPU0_RESET_N,
    output wire M_AB_CPU1_FPGA_RESET_R_N,
    input wire M_AB_CPU1_RESET_N,
    output wire M_CD_CPU0_FPGA_RESET_R_N,
    input wire M_CD_CPU0_RESET_N,
    output wire M_CD_CPU1_FPGA_RESET_R_N,
    input wire M_CD_CPU1_RESET_N,
    output wire M_EF_CPU0_FPGA_RESET_R_N,
    input wire M_EF_CPU0_RESET_N,
    output wire M_EF_CPU1_FPGA_RESET_R_N,
    input wire M_EF_CPU1_RESET_N,
    output wire M_GH_CPU0_FPGA_RESET_R_N,
    input wire M_GH_CPU0_RESET_N,
    output wire M_GH_CPU1_FPGA_RESET_R_N,
    input wire M_GH_CPU1_RESET_N,
    output wire PWRGD_CPU0_LVC1_R,
    output wire PWRGD_CPU1_LVC1_R,
    input wire PWRGD_CPUPWRGD_LVC1,
    output wire PWRGD_DRAMPWRGD_CPU0_AB_R_LVC1,
    output wire PWRGD_DRAMPWRGD_CPU0_CD_R_LVC1,
    output wire PWRGD_DRAMPWRGD_CPU0_EF_R_LVC1,
    output wire PWRGD_DRAMPWRGD_CPU0_GH_R_LVC1,
    output wire PWRGD_DRAMPWRGD_CPU1_AB_R_LVC1,
    output wire PWRGD_DRAMPWRGD_CPU1_CD_R_LVC1,
    output wire PWRGD_DRAMPWRGD_CPU1_EF_R_LVC1,
    output wire PWRGD_DRAMPWRGD_CPU1_GH_R_LVC1,
    inout wire PWRGD_FAIL_CPU0_AB_PLD,
    inout wire PWRGD_FAIL_CPU0_CD_PLD,
    inout wire PWRGD_FAIL_CPU0_EF_PLD,
    inout wire PWRGD_FAIL_CPU0_GH_PLD,
    inout wire PWRGD_FAIL_CPU1_AB_PLD,
    inout wire PWRGD_FAIL_CPU1_CD_PLD,
    inout wire PWRGD_FAIL_CPU1_EF_PLD,
    inout wire PWRGD_FAIL_CPU1_GH_PLD,
    input wire PWRGD_P1V0_BMC_AUX,
    input wire PWRGD_P1V05_PCH_AUX,
    input wire PWRGD_P1V2_BMC_AUX,
    input wire PWRGD_P1V2_MAX10_AUX_PLD_R,
    input wire PWRGD_P1V8_PCH_AUX_PLD,
    input wire PWRGD_P2V5_BMC_AUX,
    input wire PWRGD_P3V3,
    output wire PWRGD_PCH_PWROK_R,
    output wire PWRGD_PLT_AUX_CPU0_LVT3_R,
    output wire PWRGD_PLT_AUX_CPU1_LVT3_R,
    input wire PWRGD_PS_PWROK_PLD_R,
    input wire PWRGD_PVCCD_HV_CPU0,
    input wire PWRGD_PVCCD_HV_CPU1,
    input wire PWRGD_PVCCFA_EHV_CPU0,
    input wire PWRGD_PVCCFA_EHV_CPU1,
    input wire PWRGD_PVCCFA_EHV_FIVRA_CPU0,
    input wire PWRGD_PVCCFA_EHV_FIVRA_CPU1,
    input wire PWRGD_PVCCIN_CPU0,
    input wire PWRGD_PVCCIN_CPU1,
    input wire PWRGD_PVCCINFAON_CPU0,
    input wire PWRGD_PVCCINFAON_CPU1,
    input wire PWRGD_PVNN_MAIN_CPU0,
    input wire PWRGD_PVNN_MAIN_CPU1,
    input wire PWRGD_PVNN_PCH_AUX,
    input wire PWRGD_PVPP_HBM_CPU0,
    input wire PWRGD_PVPP_HBM_CPU1,
    output wire PWRGD_SYS_PWROK_R,
    output wire RST_CPU0_LVC1_R_N,
    output wire RST_CPU1_LVC1_R_N,
    input wire RST_DEDI_BUSY_PLD_N,
    output wire RST_PLD_PCIE_CPU0_DEV_PERST_N,
    output wire RST_PLD_PCIE_CPU1_DEV_PERST_N,
    output wire RST_PLD_PCIE_PCH_DEV_PERST_N,
    output wire RST_PFR_EXTRST_R_N,
    output wire RST_PFR_OVR_RTC_R,
    output wire RST_PFR_OVR_SRTC_R,
    output wire RST_PLTRST_PLD_B_N,
    input wire RST_PLTRST_PLD_N,
    output wire RST_SPI_PFR_BMC_BOOT_N,
    output wire RST_SPI_PFR_PCH_N,
    input wire SGPIO_BMC_CLK,
    output wire SGPIO_BMC_DIN_R,
    input wire SGPIO_BMC_DOUT,
    input wire SGPIO_BMC_LD_N,
    inout wire SMB_BMC_HSBP_STBY_LVC3_SCL,
    inout wire SMB_BMC_HSBP_STBY_LVC3_SDA,
    inout wire SMB_PCH_PMBUS2_STBY_LVC3_SCL,
    inout wire SMB_PCH_PMBUS2_STBY_LVC3_SDA,
    inout wire SMB_PCIE_STBY_LVC3_B_SCL,
    inout wire SMB_PCIE_STBY_LVC3_B_SDA,
    inout wire SMB_PFR_HSBP_STBY_LVC3_SCL,
    inout wire SMB_PFR_HSBP_STBY_LVC3_SDA,
    inout wire SMB_PFR_PMB1_STBY_LVC3_SCL,
    inout wire SMB_PFR_PMB1_STBY_LVC3_SDA,
    inout wire SMB_PFR_PMBUS2_STBY_LVC3_R_SCL,
    inout wire SMB_PFR_PMBUS2_STBY_LVC3_R_SDA,
    output wire SMB_PFR_RFID_STBY_LVC3_SCL,
    inout wire SMB_PFR_RFID_STBY_LVC3_SDA,
    inout wire SMB_PMBUS_SML1_STBY_LVC3_SCL,
    inout wire SMB_PMBUS_SML1_STBY_LVC3_SDA,
    input wire SMB_S3M_CPU0_SCL_LVC1,
    inout wire SMB_S3M_CPU0_SDA_LVC1,
    input wire SMB_S3M_CPU1_SCL_LVC1,
    inout wire SMB_S3M_CPU1_SDA_LVC1,
    input wire SPI_BMC_BOOT_CS_N,
    input wire SPI_BMC_BT_MUXED_MON_CLK,
    inout wire SPI_BMC_BT_MUXED_MON_IO2,
    inout wire SPI_BMC_BT_MUXED_MON_IO3,
    inout wire SPI_BMC_BT_MUXED_MON_MISO,
    inout wire SPI_BMC_BT_MUXED_MON_MOSI,
    input wire SPI_PCH_CS1_N,
    inout wire SPI_PCH_MUXED_MON_CLK,
    inout wire SPI_PCH_MUXED_MON_IO0,
    inout wire SPI_PCH_MUXED_MON_IO1,
    inout wire SPI_PCH_MUXED_MON_IO2,
    inout wire SPI_PCH_MUXED_MON_IO3,
    input wire SPI_PCH_PFR_CS0_N,
    input wire SPI_PCH_TPM_CS_N,
    inout wire SPI_PFR_BMC_BOOT_R_IO2,
    inout wire SPI_PFR_BMC_BOOT_R_IO3,
    output wire SPI_PFR_BMC_BT_SECURE_CS_R_N,
    inout wire SPI_PFR_BMC_FLASH1_BT_CLK,
    inout wire SPI_PFR_BMC_FLASH1_BT_MISO,
    inout wire SPI_PFR_BMC_FLASH1_BT_MOSI,
    inout wire SPI_PFR_PCH_R_CLK,
    inout wire SPI_PFR_PCH_R_IO0,
    inout wire SPI_PFR_PCH_R_IO1,
    inout wire SPI_PFR_PCH_R_IO2,
    inout wire SPI_PFR_PCH_R_IO3,
    output wire SPI_PFR_PCH_SECURE_CS0_R_N,
    output wire SPI_PFR_PCH_SECURE_CS1_N,
    output wire SPI_PFR_TPM_CS_R2_N,
    output wire RST_RSMRST_PLD_R_N,
    output wire RST_SRST_BMC_PLD_R_N,
    output wire FM_POSTLED_SEL,
    output wire FM_CPU_CATERR_LVT3_R_N,
    output wire FM_ADR_ACK_R,
    input wire FM_ADR_COMPLETE,
    output wire FM_ADR_TRIGGER_N,
    input wire FM_BMC_CRASHLOG_TRIG_N,
    output wire FM_PCH_CRASHLOG_TRIG_R_N,
    input wire FM_PCH_PLD_GLB_RST_WARN_N,
    input wire FM_PMBUS_ALERT_B_EN,
    input wire FM_THROTTLE_R_N,
    input wire H_CPU_CATERR_LVC1_R_N,
    output wire H_CPU_NMI_LVC1_R,
    input wire IRQ_BMC_CPU_NMI,
    input wire IRQ_PCH_CPU_NMI_EVENT_N,
    inout wire IRQ_SML1_PMBUS_PLD_ALERT_N,
    output wire FM_CPU1_DIMM_CH1_4_FAULT_LED_SEL,
    output wire FM_CPU1_DIMM_CH5_8_FAULT_LED_SEL,
    output wire FM_CPU0_DIMM_CH1_4_FAULT_LED_SEL,
    output wire FM_CPU0_DIMM_CH5_8_FAULT_LED_SEL,
    output wire FM_POST_7SEG1_SEL_N,
    output wire FM_POST_7SEG2_SEL_N,
    output wire FM_FAN_FAULT_LED_SEL_R_N,
    input wire H_CPU_ERR0_LVC1_R_N,
    input wire H_CPU_ERR1_LVC1_R_N,
    input wire H_CPU_ERR2_LVC1_R_N,
    output wire FM_CPU_ERR0_LVT3_N,
    output wire FM_CPU_ERR1_LVT3_N,
    output wire FM_CPU_ERR2_LVT3_N,
    input wire FM_DIS_PS_PWROK_DLY,
    output wire FM_HBM2_HBM3_VPP_SEL,
    output wire PWRGD_S0_PWROK_CPU0_LVC1_R,
    output wire PWRGD_S0_PWROK_CPU1_LVC1_R,
    input wire SGPIO_DEBUG_PLD_CLK,
    input wire SGPIO_DEBUG_PLD_DOUT,
    input wire SGPIO_DEBUG_PLD_LD,
    output wire SGPIO_DEBUG_PLD_DIN,
    input wire FP_BMC_PWR_BTN_R2_N,
    input wire FM_VAL_BOARD_PRSNT_N,
    input wire FM_ADR_MODE0,
    input wire FM_ADR_MODE1,
    output wire IRQ_BMC_PCH_NMI,
    input wire FM_S3M_CPU0_CPLD_CRC_ERROR,
    input wire FM_S3M_CPU1_CPLD_CRC_ERROR,
    input wire SGPIO_IDV_CLK_R,
    input wire SGPIO_IDV_DOUT_R,
    output wire SGPIO_IDV_DIN_R,
    input wire SGPIO_IDV_LD_R_N

);

    // Clocks and resets
    wire pll_locked;
    wire clk2M;
    wire clk50M;
    wire sys_clk;
    wire spi_clk;
    wire clk2M_reset_sync_n;
    wire clk50M_reset_sync_n;
    wire sys_clk_reset_sync_n;
    wire spi_clk_reset_sync_n;
    
    // BMC/PCH reset generation signals from common core
    wire wRST_RSMRST_PLD_R_N_REQ;
    wire wRST_SRST_BMC_PLD_R_N_REQ;
   
    // LED Control from common core
    wire wLED_CONTROL_0;
    wire wLED_CONTROL_1;
    wire wLED_CONTROL_2;
    wire wLED_CONTROL_3;
    wire wLED_CONTROL_4;
    wire wLED_CONTROL_5;
    wire wLED_CONTROL_6;
    wire wLED_CONTROL_7;
    wire wFM_POST_7SEG1_SEL_N;
    wire wFM_POST_7SEG2_SEL_N;
    wire wFM_POSTLED_SEL;

    // HPFR signals from the common core
    // TODO Connect to common core when changes have been made
    wire wHPFR_IN;
    wire wHPFR_OUT;
    wire wLEGACY;
    wire wHPFR_ACTIVE;
    wire wRST_PLTRST_PLD_N;

    // Clocks and reset generator
    pfr_sys_clocks_reset u_pfr_sys_clocks_reset (
        .refclk(CLK_25M_OSC_MAIN_FPGA),
        .pll_reset(!PWRGD_P1V2_MAX10_AUX_PLD_R),
        .pll_locked(pll_locked),
        .clk2M(clk2M),
        .clk50M(clk50M),
        .sys_clk(sys_clk),
        .spi_clk(spi_clk),
        .clk2M_reset_sync_n(clk2M_reset_sync_n),
        .clk50M_reset_sync_n(clk50M_reset_sync_n),
        .sys_clk_reset_sync_n(sys_clk_reset_sync_n),
        .spi_clk_reset_sync_n(spi_clk_reset_sync_n)
    );
        
    // Instantiate the common core
    Archer_City_Main_wrapper u_common_core (
        .iClk_2M(clk2M),
        .iClk_50M(clk50M),
        .ipll_locked(pll_locked),
        
        .RST_RSMRST_PLD_R_N(RST_RSMRST_PLD_R_N),
        .RST_SRST_BMC_PLD_R_N(RST_SRST_BMC_PLD_R_N),
        .RST_RSMRST_PLD_R_N_REQ(wRST_RSMRST_PLD_R_N_REQ),
        .RST_SRST_BMC_PLD_R_N_REQ(wRST_SRST_BMC_PLD_R_N_REQ),
        .RST_PLTRST_PLD_N(wRST_PLTRST_PLD_N),
        
        .LED_CONTROL_0(wLED_CONTROL_0),
        .LED_CONTROL_1(wLED_CONTROL_1),
        .LED_CONTROL_2(wLED_CONTROL_2),
        .LED_CONTROL_3(wLED_CONTROL_3),
        .LED_CONTROL_4(wLED_CONTROL_4),
        .LED_CONTROL_5(wLED_CONTROL_5),
        .LED_CONTROL_6(wLED_CONTROL_6),
        .LED_CONTROL_7(wLED_CONTROL_7),
        .FM_POST_7SEG1_SEL_N(wFM_POST_7SEG1_SEL_N),
        .FM_POST_7SEG2_SEL_N(wFM_POST_7SEG2_SEL_N),
        .FM_POSTLED_SEL(wFM_POSTLED_SEL),
        .HPFR_TO_MISC(wHPFR_OUT),
        .HPFR_FROM_MISC(wHPFR_IN),
        .FM_MODULAR_LEGACY(wLEGACY),
        .FM_MODULAR_STANDALONE(wHPFR_ACTIVE),
        
        .FM_AUX_SW_EN(FM_AUX_SW_EN),
        .FM_BMC_NMI_PCH_EN(FM_BMC_NMI_PCH_EN),
        .FM_BMC_ONCTL_N_PLD(FM_BMC_ONCTL_N_PLD),
        .FM_BMC_PFR_PWRBTN_OUT_R_N(FM_BMC_PFR_PWRBTN_OUT_R_N),
        .FM_BMC_PWRBTN_OUT_N(FM_BMC_PWRBTN_OUT_N),
        .FM_CPU0_INTR_PRSNT(FM_CPU0_INTR_PRSNT),
        .FM_CPU0_PKGID0(FM_CPU0_PKGID0),
        .FM_CPU0_PKGID1(FM_CPU0_PKGID1),
        .FM_CPU0_PKGID2(FM_CPU0_PKGID2),
        .FM_CPU0_PROC_ID0(FM_CPU0_PROC_ID0),
        .FM_CPU0_PROC_ID1(FM_CPU0_PROC_ID1),
        .FM_CPU0_SKTOCC_LVT3_PLD_N(FM_CPU0_SKTOCC_LVT3_PLD_N),
        .FM_CPU1_PKGID0(FM_CPU1_PKGID0),
        .FM_CPU1_PKGID1(FM_CPU1_PKGID1),
        .FM_CPU1_PKGID2(FM_CPU1_PKGID2),
        .FM_CPU1_PROC_ID0(FM_CPU1_PROC_ID0),
        .FM_CPU1_PROC_ID1(FM_CPU1_PROC_ID1),
        .FM_CPU1_SKTOCC_LVT3_PLD_N(FM_CPU1_SKTOCC_LVT3_PLD_N),
        .FM_DIMM_12V_CPS_S5_N(FM_DIMM_12V_CPS_S5_N),
        .FM_FORCE_PWRON_LVC3(FM_FORCE_PWRON_LVC3),
        .FM_P1V0_BMC_AUX_EN(FM_P1V0_BMC_AUX_EN),
        .FM_P1V05_PCH_AUX_EN(FM_P1V05_PCH_AUX_EN),
        .FM_P1V2_BMC_AUX_EN(FM_P1V2_BMC_AUX_EN),
        .FM_P2V5_BMC_AUX_EN(FM_P2V5_BMC_AUX_EN),
        .FM_P5V_EN(FM_P5V_EN),
        .FM_PCH_P1V8_AUX_EN(FM_PCH_P1V8_AUX_EN),
        .FM_PCH_PRSNT_N(FM_PCH_PRSNT_N),
        .FM_PFR_MUX_OE_CTL_PLD(FM_PFR_MUX_OE_CTL_PLD),
        .FM_PLD_CLK_25M_R_EN(FM_PLD_CLK_25M_R_EN),
        .FM_PLD_CLKS_DEV_R_EN(FM_PLD_CLKS_DEV_R_EN),
        .FM_PLD_HEARTBEAT_LVC3(FM_PLD_HEARTBEAT_LVC3),
        .FM_PLD_REV_N(FM_PLD_REV_N),
        .FM_PS_EN_PLD_R(FM_PS_EN_PLD_R),
        .FM_PVCCD_HV_CPU0_EN(FM_PVCCD_HV_CPU0_EN),
        .FM_PVCCD_HV_CPU1_EN(FM_PVCCD_HV_CPU1_EN),
        .FM_PVCCFA_EHV_CPU0_R_EN(FM_PVCCFA_EHV_CPU0_R_EN),
        .FM_PVCCFA_EHV_CPU1_R_EN(FM_PVCCFA_EHV_CPU1_R_EN),
        .FM_PVCCFA_EHV_FIVRA_CPU0_R_EN(FM_PVCCFA_EHV_FIVRA_CPU0_R_EN),
        .FM_PVCCFA_EHV_FIVRA_CPU1_R_EN(FM_PVCCFA_EHV_FIVRA_CPU1_R_EN),
        .FM_PVCCIN_CPU0_R_EN(FM_PVCCIN_CPU0_R_EN),
        .FM_PVCCIN_CPU1_R_EN(FM_PVCCIN_CPU1_R_EN),
        .FM_PVCCINFAON_CPU0_R_EN(FM_PVCCINFAON_CPU0_R_EN),
        .FM_PVCCINFAON_CPU1_R_EN(FM_PVCCINFAON_CPU1_R_EN),
        .FM_PVNN_MAIN_CPU0_EN(FM_PVNN_MAIN_CPU0_EN),
        .FM_PVNN_MAIN_CPU1_EN(FM_PVNN_MAIN_CPU1_EN),
        .FM_PVNN_PCH_AUX_EN(FM_PVNN_PCH_AUX_EN),
        .FM_PVPP_HBM_CPU0_EN(FM_PVPP_HBM_CPU0_EN),
        .FM_PVPP_HBM_CPU1_EN(FM_PVPP_HBM_CPU1_EN),
        .FM_RST_PERST_BIT0(FM_RST_PERST_BIT0),
        .FM_RST_PERST_BIT1(FM_RST_PERST_BIT1),
        .FM_RST_PERST_BIT2(FM_RST_PERST_BIT2),
        .FM_SLP_SUS_RSM_RST_N(FM_SLP_SUS_RSM_RST_N),
        .FM_SLPS3_PLD_N(FM_SLPS3_PLD_N),
        .FM_SLPS4_PLD_N(FM_SLPS4_PLD_N),
        .FM_SX_SW_P12V_R_EN(FM_SX_SW_P12V_R_EN),
        .FM_SX_SW_P12V_STBY_R_EN(FM_SX_SW_P12V_STBY_R_EN),
        .FM_SYS_THROTTLE_R_N(FM_SYS_THROTTLE_R_N),
        .FM_THERMTRIP_DLY_LVC1_R_N(FM_THERMTRIP_DLY_LVC1_R_N),
        .H_CPU0_MEMHOT_IN_LVC1_R_N(H_CPU0_MEMHOT_IN_LVC1_R_N),
        .H_CPU0_MEMHOT_OUT_LVC1_N(H_CPU0_MEMHOT_OUT_LVC1_N),
        .H_CPU0_MEMTRIP_LVC1_N(H_CPU0_MEMTRIP_LVC1_N),
        .H_CPU0_MON_FAIL_PLD_LVC1_N(H_CPU0_MON_FAIL_PLD_LVC1_N),
        .H_CPU0_PROCHOT_LVC1_R_N(H_CPU0_PROCHOT_LVC1_R_N),
        .H_CPU0_THERMTRIP_LVC1_N(H_CPU0_THERMTRIP_LVC1_N),
        .H_CPU1_MEMHOT_IN_LVC1_R_N(H_CPU1_MEMHOT_IN_LVC1_R_N),
        .H_CPU1_MEMHOT_OUT_LVC1_N(H_CPU1_MEMHOT_OUT_LVC1_N),
        .H_CPU1_MEMTRIP_LVC1_N(H_CPU1_MEMTRIP_LVC1_N),
        .H_CPU1_MON_FAIL_PLD_LVC1_N(H_CPU1_MON_FAIL_PLD_LVC1_N),
        .H_CPU1_PROCHOT_LVC1_R_N(H_CPU1_PROCHOT_LVC1_R_N),
        .H_CPU1_THERMTRIP_LVC1_N(H_CPU1_THERMTRIP_LVC1_N),
        .IRQ_CPU0_MEM_VRHOT_N(IRQ_CPU0_MEM_VRHOT_N),
        .IRQ_CPU0_VRHOT_N(IRQ_CPU0_VRHOT_N),
        .IRQ_CPU1_MEM_VRHOT_N(IRQ_CPU1_MEM_VRHOT_N),
        .IRQ_CPU1_VRHOT_N(IRQ_CPU1_VRHOT_N),
        .M_AB_CPU0_FPGA_RESET_R_N(M_AB_CPU0_FPGA_RESET_R_N),
        .M_AB_CPU0_RESET_N(M_AB_CPU0_RESET_N),
        .M_AB_CPU1_FPGA_RESET_R_N(M_AB_CPU1_FPGA_RESET_R_N),
        .M_AB_CPU1_RESET_N(M_AB_CPU1_RESET_N),
        .M_CD_CPU0_FPGA_RESET_R_N(M_CD_CPU0_FPGA_RESET_R_N),
        .M_CD_CPU0_RESET_N(M_CD_CPU0_RESET_N),
        .M_CD_CPU1_FPGA_RESET_R_N(M_CD_CPU1_FPGA_RESET_R_N),
        .M_CD_CPU1_RESET_N(M_CD_CPU1_RESET_N),
        .M_EF_CPU0_FPGA_RESET_R_N(M_EF_CPU0_FPGA_RESET_R_N),
        .M_EF_CPU0_RESET_N(M_EF_CPU0_RESET_N),
        .M_EF_CPU1_FPGA_RESET_R_N(M_EF_CPU1_FPGA_RESET_R_N),
        .M_EF_CPU1_RESET_N(M_EF_CPU1_RESET_N),
        .M_GH_CPU0_FPGA_RESET_R_N(M_GH_CPU0_FPGA_RESET_R_N),
        .M_GH_CPU0_RESET_N(M_GH_CPU0_RESET_N),
        .M_GH_CPU1_FPGA_RESET_R_N(M_GH_CPU1_FPGA_RESET_R_N),
        .M_GH_CPU1_RESET_N(M_GH_CPU1_RESET_N),
        .PWRGD_CPU0_LVC1_R(PWRGD_CPU0_LVC1_R),
        .PWRGD_CPU1_LVC1_R(PWRGD_CPU1_LVC1_R),
        .PWRGD_CPUPWRGD_LVC1(PWRGD_CPUPWRGD_LVC1),
        .PWRGD_DRAMPWRGD_CPU0_AB_R_LVC1(PWRGD_DRAMPWRGD_CPU0_AB_R_LVC1),
        .PWRGD_DRAMPWRGD_CPU0_CD_R_LVC1(PWRGD_DRAMPWRGD_CPU0_CD_R_LVC1),
        .PWRGD_DRAMPWRGD_CPU0_EF_R_LVC1(PWRGD_DRAMPWRGD_CPU0_EF_R_LVC1),
        .PWRGD_DRAMPWRGD_CPU0_GH_R_LVC1(PWRGD_DRAMPWRGD_CPU0_GH_R_LVC1),
        .PWRGD_DRAMPWRGD_CPU1_AB_R_LVC1(PWRGD_DRAMPWRGD_CPU1_AB_R_LVC1),
        .PWRGD_DRAMPWRGD_CPU1_CD_R_LVC1(PWRGD_DRAMPWRGD_CPU1_CD_R_LVC1),
        .PWRGD_DRAMPWRGD_CPU1_EF_R_LVC1(PWRGD_DRAMPWRGD_CPU1_EF_R_LVC1),
        .PWRGD_DRAMPWRGD_CPU1_GH_R_LVC1(PWRGD_DRAMPWRGD_CPU1_GH_R_LVC1),
        .PWRGD_FAIL_CPU0_AB_PLD(PWRGD_FAIL_CPU0_AB_PLD),
        .PWRGD_FAIL_CPU0_CD_PLD(PWRGD_FAIL_CPU0_CD_PLD),
        .PWRGD_FAIL_CPU0_EF_PLD(PWRGD_FAIL_CPU0_EF_PLD),
        .PWRGD_FAIL_CPU0_GH_PLD(PWRGD_FAIL_CPU0_GH_PLD),
        .PWRGD_FAIL_CPU1_AB_PLD(PWRGD_FAIL_CPU1_AB_PLD),
        .PWRGD_FAIL_CPU1_CD_PLD(PWRGD_FAIL_CPU1_CD_PLD),
        .PWRGD_FAIL_CPU1_EF_PLD(PWRGD_FAIL_CPU1_EF_PLD),
        .PWRGD_FAIL_CPU1_GH_PLD(PWRGD_FAIL_CPU1_GH_PLD),
        .PWRGD_P1V0_BMC_AUX(PWRGD_P1V0_BMC_AUX),
        .PWRGD_P1V05_PCH_AUX(PWRGD_P1V05_PCH_AUX),
        .PWRGD_P1V2_BMC_AUX(PWRGD_P1V2_BMC_AUX),
        .PWRGD_P1V2_MAX10_AUX_PLD_R(PWRGD_P1V2_MAX10_AUX_PLD_R),
        .PWRGD_P1V8_PCH_AUX_PLD(PWRGD_P1V8_PCH_AUX_PLD),
        .PWRGD_P2V5_BMC_AUX(PWRGD_P2V5_BMC_AUX),
        .PWRGD_P3V3(PWRGD_P3V3),
        .PWRGD_PCH_PWROK_R(PWRGD_PCH_PWROK_R),
        .PWRGD_PLT_AUX_CPU0_LVT3_R(PWRGD_PLT_AUX_CPU0_LVT3_R),
        .PWRGD_PLT_AUX_CPU1_LVT3_R(PWRGD_PLT_AUX_CPU1_LVT3_R),
        .PWRGD_PS_PWROK_PLD_R(PWRGD_PS_PWROK_PLD_R),
        .PWRGD_PVCCD_HV_CPU0(PWRGD_PVCCD_HV_CPU0),
        .PWRGD_PVCCD_HV_CPU1(PWRGD_PVCCD_HV_CPU1),
        .PWRGD_PVCCFA_EHV_CPU0(PWRGD_PVCCFA_EHV_CPU0),
        .PWRGD_PVCCFA_EHV_CPU1(PWRGD_PVCCFA_EHV_CPU1),
        .PWRGD_PVCCFA_EHV_FIVRA_CPU0(PWRGD_PVCCFA_EHV_FIVRA_CPU0),
        .PWRGD_PVCCFA_EHV_FIVRA_CPU1(PWRGD_PVCCFA_EHV_FIVRA_CPU1),
        .PWRGD_PVCCIN_CPU0(PWRGD_PVCCIN_CPU0),
        .PWRGD_PVCCIN_CPU1(PWRGD_PVCCIN_CPU1),
        .PWRGD_PVCCINFAON_CPU0(PWRGD_PVCCINFAON_CPU0),
        .PWRGD_PVCCINFAON_CPU1(PWRGD_PVCCINFAON_CPU1),
        .PWRGD_PVNN_MAIN_CPU0(PWRGD_PVNN_MAIN_CPU0),
        .PWRGD_PVNN_MAIN_CPU1(PWRGD_PVNN_MAIN_CPU1),
        .PWRGD_PVNN_PCH_AUX(PWRGD_PVNN_PCH_AUX),
        .PWRGD_PVPP_HBM_CPU0(PWRGD_PVPP_HBM_CPU0),
        .PWRGD_PVPP_HBM_CPU1(PWRGD_PVPP_HBM_CPU1),
        .PWRGD_SYS_PWROK_R(PWRGD_SYS_PWROK_R),
        .RST_CPU0_LVC1_R_N(RST_CPU0_LVC1_R_N),
        .RST_CPU1_LVC1_R_N(RST_CPU1_LVC1_R_N),
        .RST_DEDI_BUSY_PLD_N(RST_DEDI_BUSY_PLD_N),
        .RST_PLD_PCIE_CPU0_DEV_PERST_N(RST_PLD_PCIE_CPU0_DEV_PERST_N),
        .RST_PLD_PCIE_CPU1_DEV_PERST_N(RST_PLD_PCIE_CPU1_DEV_PERST_N),
        .RST_PLD_PCIE_PCH_DEV_PERST_N(RST_PLD_PCIE_PCH_DEV_PERST_N),
        .RST_PLTRST_PLD_B_N(RST_PLTRST_PLD_B_N),
        .SGPIO_BMC_CLK(SGPIO_BMC_CLK),
        .SGPIO_BMC_DIN_R(SGPIO_BMC_DIN_R),
        .SGPIO_BMC_DOUT(SGPIO_BMC_DOUT),
        .SGPIO_BMC_LD_N(SGPIO_BMC_LD_N),
        .SMB_S3M_CPU0_SCL_LVC1(SMB_S3M_CPU0_SCL_LVC1),
        .SMB_S3M_CPU0_SDA_LVC1(SMB_S3M_CPU0_SDA_LVC1),
        .SMB_S3M_CPU1_SCL_LVC1(SMB_S3M_CPU1_SCL_LVC1),
        .SMB_S3M_CPU1_SDA_LVC1(SMB_S3M_CPU1_SDA_LVC1),
        .FM_CPU_CATERR_LVT3_R_N(FM_CPU_CATERR_LVT3_R_N),
        .FM_ADR_ACK_R(FM_ADR_ACK_R),
        .FM_ADR_COMPLETE(FM_ADR_COMPLETE),
        .FM_ADR_TRIGGER_N(FM_ADR_TRIGGER_N),
        .FM_BMC_CRASHLOG_TRIG_N(FM_BMC_CRASHLOG_TRIG_N),
        .FM_PCH_CRASHLOG_TRIG_R_N(FM_PCH_CRASHLOG_TRIG_R_N),
        .FM_PCH_PLD_GLB_RST_WARN_N(FM_PCH_PLD_GLB_RST_WARN_N),
        .FM_PMBUS_ALERT_B_EN(FM_PMBUS_ALERT_B_EN),
        .FM_THROTTLE_R_N(FM_THROTTLE_R_N),
        .H_CPU_CATERR_LVC1_R_N(H_CPU_CATERR_LVC1_R_N),
        .H_CPU_NMI_LVC1_R(H_CPU_NMI_LVC1_R),
        .IRQ_BMC_CPU_NMI(IRQ_BMC_CPU_NMI),
        .IRQ_PCH_CPU_NMI_EVENT_N(IRQ_PCH_CPU_NMI_EVENT_N),
        .IRQ_SML1_PMBUS_PLD_ALERT_N(IRQ_SML1_PMBUS_PLD_ALERT_N),
        .FM_CPU1_DIMM_CH1_4_FAULT_LED_SEL(FM_CPU1_DIMM_CH1_4_FAULT_LED_SEL),
        .FM_CPU1_DIMM_CH5_8_FAULT_LED_SEL(FM_CPU1_DIMM_CH5_8_FAULT_LED_SEL),
        .FM_CPU0_DIMM_CH1_4_FAULT_LED_SEL(FM_CPU0_DIMM_CH1_4_FAULT_LED_SEL),
        .FM_CPU0_DIMM_CH5_8_FAULT_LED_SEL(FM_CPU0_DIMM_CH5_8_FAULT_LED_SEL),
        .FM_FAN_FAULT_LED_SEL_R_N(FM_FAN_FAULT_LED_SEL_R_N),
        .H_CPU_ERR0_LVC1_R_N(H_CPU_ERR0_LVC1_R_N),
        .H_CPU_ERR1_LVC1_R_N(H_CPU_ERR1_LVC1_R_N),
        .H_CPU_ERR2_LVC1_R_N(H_CPU_ERR2_LVC1_R_N),
        .FM_CPU_ERR0_LVT3_N(FM_CPU_ERR0_LVT3_N),
        .FM_CPU_ERR1_LVT3_N(FM_CPU_ERR1_LVT3_N),
        .FM_CPU_ERR2_LVT3_N(FM_CPU_ERR2_LVT3_N),
        .FM_DIS_PS_PWROK_DLY(FM_DIS_PS_PWROK_DLY),
        .FM_HBM2_HBM3_VPP_SEL(FM_HBM2_HBM3_VPP_SEL),
        .PWRGD_S0_PWROK_CPU0_LVC1_R(PWRGD_S0_PWROK_CPU0_LVC1_R),
        .PWRGD_S0_PWROK_CPU1_LVC1_R(PWRGD_S0_PWROK_CPU1_LVC1_R),
        .SGPIO_DEBUG_PLD_CLK(SGPIO_DEBUG_PLD_CLK),
        .SGPIO_DEBUG_PLD_DOUT(SGPIO_DEBUG_PLD_DOUT),
        .SGPIO_DEBUG_PLD_LD(SGPIO_DEBUG_PLD_LD),
        .SGPIO_DEBUG_PLD_DIN(SGPIO_DEBUG_PLD_DIN),
        .FP_BMC_PWR_BTN_R2_N(FP_BMC_PWR_BTN_R2_N),
        .FM_VAL_BOARD_PRSNT_N(FM_VAL_BOARD_PRSNT_N),
        .FM_ADR_MODE0(FM_ADR_MODE0),
        .FM_ADR_MODE1(FM_ADR_MODE1),
        .IRQ_BMC_PCH_NMI(IRQ_BMC_PCH_NMI),
        .FM_S3M_CPU0_CPLD_CRC_ERROR(FM_S3M_CPU0_CPLD_CRC_ERROR),
        .FM_S3M_CPU1_CPLD_CRC_ERROR(FM_S3M_CPU1_CPLD_CRC_ERROR),
        .SGPIO_IDV_CLK_R(SGPIO_IDV_CLK_R),
        .SGPIO_IDV_DOUT_R(SGPIO_IDV_DOUT_R),
        .SGPIO_IDV_DIN_R(SGPIO_IDV_DIN_R),
        .SGPIO_IDV_LD_R_N(SGPIO_IDV_LD_R_N)

    );

    recovery_core u_core (

        .clk2M(clk2M),
        .clk50M(clk50M),
        .sys_clk(sys_clk),
        .spi_clk(spi_clk),
        .clk2M_reset_sync_n(clk2M_reset_sync_n),
        .clk50M_reset_sync_n(clk50M_reset_sync_n),
        .sys_clk_reset_sync_n(sys_clk_reset_sync_n),
        .spi_clk_reset_sync_n(spi_clk_reset_sync_n),
        
        .cc_RST_RSMRST_PLD_R_N(wRST_RSMRST_PLD_R_N_REQ),
        .cc_RST_SRST_BMC_PLD_R_N(wRST_SRST_BMC_PLD_R_N_REQ),
        .cc_RST_PLTRST_PLD_N(wRST_PLTRST_PLD_N),
        
        .ccLED_CONTROL_0(wLED_CONTROL_0),
        .ccLED_CONTROL_1(wLED_CONTROL_1),
        .ccLED_CONTROL_2(wLED_CONTROL_2),
        .ccLED_CONTROL_3(wLED_CONTROL_3),
        .ccLED_CONTROL_4(wLED_CONTROL_4),
        .ccLED_CONTROL_5(wLED_CONTROL_5),
        .ccLED_CONTROL_6(wLED_CONTROL_6),
        .ccLED_CONTROL_7(wLED_CONTROL_7),
        .ccFM_POST_7SEG1_SEL_N(wFM_POST_7SEG1_SEL_N),
        .ccFM_POST_7SEG2_SEL_N(wFM_POST_7SEG2_SEL_N),
        .ccFM_POSTLED_SEL(wFM_POSTLED_SEL),

        .ccHPFR_IN(wHPFR_IN),
        .ccHPFR_OUT(wHPFR_OUT),
        .ccLEGACY(wLEGACY),
        .ccHPFR_ACTIVE(wHPFR_ACTIVE),


        .FAN_BMC_PWM_R(FAN_BMC_PWM_R),
        .FM_ME_AUTHN_FAIL(FM_ME_AUTHN_FAIL),
        .FM_ME_BT_DONE(FM_ME_BT_DONE),
        .FM_PFR_DSW_PWROK_N(FM_PFR_DSW_PWROK_N),
        .FM_PFR_FORCE_RECOVERY_N(FM_PFR_FORCE_RECOVERY_N),
        .FM_PFR_ON_R(FM_PFR_ON_R),
        .FM_PFR_POSTCODE_SEL_N(FM_PFR_POSTCODE_SEL_N),
        .FM_PFR_RNDGEN_AUX(FM_PFR_RNDGEN_AUX),
        .FM_PFR_SLP_SUS_EN_R_N(FM_PFR_SLP_SUS_EN_R_N),
        .FM_PFR_TM1_HOLD_N(FM_PFR_TM1_HOLD_N),
        .FM_SPI_PFR_BMC_BT_MASTER_SEL_R(FM_SPI_PFR_BMC_BT_MASTER_SEL_R),
        .FM_SPI_PFR_PCH_MASTER_SEL_R(FM_SPI_PFR_PCH_MASTER_SEL_R),
        .FP_ID_LED_N(FP_ID_LED_N),
        .FP_ID_LED_PFR_N(FP_ID_LED_PFR_N),
        .FP_LED_STATUS_AMBER_N(FP_LED_STATUS_AMBER_N),
        .FP_LED_STATUS_AMBER_PFR_N(FP_LED_STATUS_AMBER_PFR_N),
        .FP_LED_STATUS_GREEN_N(FP_LED_STATUS_GREEN_N),
        .FP_LED_STATUS_GREEN_PFR_N(FP_LED_STATUS_GREEN_PFR_N),
        .LED_CONTROL_0(LED_CONTROL_0),
        .LED_CONTROL_1(LED_CONTROL_1),
        .LED_CONTROL_2(LED_CONTROL_2),
        .LED_CONTROL_3(LED_CONTROL_3),
        .LED_CONTROL_4(LED_CONTROL_4),
        .LED_CONTROL_5(LED_CONTROL_5),
        .LED_CONTROL_6(LED_CONTROL_6),
        .LED_CONTROL_7(LED_CONTROL_7),
        .RST_PFR_EXTRST_R_N(RST_PFR_EXTRST_R_N),
        .RST_PFR_OVR_RTC_R(RST_PFR_OVR_RTC_R),
        .RST_PFR_OVR_SRTC_R(RST_PFR_OVR_SRTC_R),
        .RST_PLTRST_PLD_N(RST_PLTRST_PLD_N),
        .RST_SPI_PFR_BMC_BOOT_N(RST_SPI_PFR_BMC_BOOT_N),
        .RST_SPI_PFR_PCH_N(RST_SPI_PFR_PCH_N),
        .SMB_BMC_HSBP_STBY_LVC3_SCL(SMB_BMC_HSBP_STBY_LVC3_SCL),
        .SMB_BMC_HSBP_STBY_LVC3_SDA(SMB_BMC_HSBP_STBY_LVC3_SDA),
        .SMB_PCH_PMBUS2_STBY_LVC3_SCL(SMB_PCH_PMBUS2_STBY_LVC3_SCL),
        .SMB_PCH_PMBUS2_STBY_LVC3_SDA(SMB_PCH_PMBUS2_STBY_LVC3_SDA),
        .SMB_PCIE_STBY_LVC3_B_SCL(SMB_PCIE_STBY_LVC3_B_SCL),
        .SMB_PCIE_STBY_LVC3_B_SDA(SMB_PCIE_STBY_LVC3_B_SDA),
        .SMB_PFR_HSBP_STBY_LVC3_SCL(SMB_PFR_HSBP_STBY_LVC3_SCL),
        .SMB_PFR_HSBP_STBY_LVC3_SDA(SMB_PFR_HSBP_STBY_LVC3_SDA),
        .SMB_PFR_PMB1_STBY_LVC3_SCL(SMB_PFR_PMB1_STBY_LVC3_SCL),
        .SMB_PFR_PMB1_STBY_LVC3_SDA(SMB_PFR_PMB1_STBY_LVC3_SDA),
        .SMB_PFR_PMBUS2_STBY_LVC3_R_SCL(SMB_PFR_PMBUS2_STBY_LVC3_R_SCL),
        .SMB_PFR_PMBUS2_STBY_LVC3_R_SDA(SMB_PFR_PMBUS2_STBY_LVC3_R_SDA),
        .SMB_PFR_RFID_STBY_LVC3_SCL(SMB_PFR_RFID_STBY_LVC3_SCL),
        .SMB_PFR_RFID_STBY_LVC3_SDA(SMB_PFR_RFID_STBY_LVC3_SDA),
        .SMB_PMBUS_SML1_STBY_LVC3_SCL(SMB_PMBUS_SML1_STBY_LVC3_SCL),
        .SMB_PMBUS_SML1_STBY_LVC3_SDA(SMB_PMBUS_SML1_STBY_LVC3_SDA),
        .SMB_S3M_CPU0_SCL_LVC1(SMB_S3M_CPU0_SCL_LVC1),
        .SMB_S3M_CPU0_SDA_LVC1(SMB_S3M_CPU0_SDA_LVC1),
        .SPI_BMC_BOOT_CS_N(SPI_BMC_BOOT_CS_N),
        .SPI_BMC_BT_MUXED_MON_CLK(SPI_BMC_BT_MUXED_MON_CLK),
        .SPI_BMC_BT_MUXED_MON_IO2(SPI_BMC_BT_MUXED_MON_IO2),
        .SPI_BMC_BT_MUXED_MON_IO3(SPI_BMC_BT_MUXED_MON_IO3),
        .SPI_BMC_BT_MUXED_MON_MISO(SPI_BMC_BT_MUXED_MON_MISO),
        .SPI_BMC_BT_MUXED_MON_MOSI(SPI_BMC_BT_MUXED_MON_MOSI),
        .SPI_PCH_CS1_N(SPI_PCH_CS1_N),
        .SPI_PCH_MUXED_MON_CLK(SPI_PCH_MUXED_MON_CLK),
        .SPI_PCH_MUXED_MON_IO0(SPI_PCH_MUXED_MON_IO0),
        .SPI_PCH_MUXED_MON_IO1(SPI_PCH_MUXED_MON_IO1),
        .SPI_PCH_MUXED_MON_IO2(SPI_PCH_MUXED_MON_IO2),
        .SPI_PCH_MUXED_MON_IO3(SPI_PCH_MUXED_MON_IO3),
        .SPI_PCH_PFR_CS0_N(SPI_PCH_PFR_CS0_N),
        .SPI_PCH_TPM_CS_N(SPI_PCH_TPM_CS_N),
        .SPI_PFR_BMC_BOOT_R_IO2(SPI_PFR_BMC_BOOT_R_IO2),
        .SPI_PFR_BMC_BOOT_R_IO3(SPI_PFR_BMC_BOOT_R_IO3),
        .SPI_PFR_BMC_BT_SECURE_CS_R_N(SPI_PFR_BMC_BT_SECURE_CS_R_N),
        .SPI_PFR_BMC_FLASH1_BT_CLK(SPI_PFR_BMC_FLASH1_BT_CLK),
        .SPI_PFR_BMC_FLASH1_BT_MISO(SPI_PFR_BMC_FLASH1_BT_MISO),
        .SPI_PFR_BMC_FLASH1_BT_MOSI(SPI_PFR_BMC_FLASH1_BT_MOSI),
        .SPI_PFR_PCH_R_CLK(SPI_PFR_PCH_R_CLK),
        .SPI_PFR_PCH_R_IO0(SPI_PFR_PCH_R_IO0),
        .SPI_PFR_PCH_R_IO1(SPI_PFR_PCH_R_IO1),
        .SPI_PFR_PCH_R_IO2(SPI_PFR_PCH_R_IO2),
        .SPI_PFR_PCH_R_IO3(SPI_PFR_PCH_R_IO3),
        .SPI_PFR_PCH_SECURE_CS0_R_N(SPI_PFR_PCH_SECURE_CS0_R_N),
        .SPI_PFR_PCH_SECURE_CS1_N(SPI_PFR_PCH_SECURE_CS1_N),
        .SPI_PFR_TPM_CS_R2_N(SPI_PFR_TPM_CS_R2_N),
        .RST_RSMRST_PLD_R_N(RST_RSMRST_PLD_R_N),
        .RST_SRST_BMC_PLD_R_N(RST_SRST_BMC_PLD_R_N),
        .FM_POSTLED_SEL(FM_POSTLED_SEL),
        .FM_POST_7SEG1_SEL_N(FM_POST_7SEG1_SEL_N),
        .FM_POST_7SEG2_SEL_N(FM_POST_7SEG2_SEL_N)

    );



endmodule
