`timescale 1 ps / 1 ps
`default_nettype none

module pfr_core (
    input wire clk2M,
    input wire clk50M,
    input wire sys_clk,
    input wire clk2M_reset_sync_n,
    input wire clk50M_reset_sync_n,
    input wire sys_clk_reset_sync_n,

    input wire cc_RST_RSMRST_PLD_R_N,
    input wire cc_RST_SRST_BMC_PLD_R_N,
    output wire cc_RST_PLTRST_PLD_N,

    input wire i1mSCE,
    input wire i1SCE,

    input wire ccLED_CONTROL_0,
    input wire ccLED_CONTROL_1,
    input wire ccLED_CONTROL_2,
    input wire ccLED_CONTROL_3,
    input wire ccLED_CONTROL_4,
    input wire ccLED_CONTROL_5,
    input wire ccLED_CONTROL_6,
    input wire ccLED_CONTROL_7,
    input wire ccFM_POST_7SEG1_SEL_N,
    input wire ccFM_POST_7SEG2_SEL_N,
    input wire ccFM_POSTLED_SEL,
    
    output wire FAN_BMC_PWM_R,
    input wire FM_ME_AUTHN_FAIL,
    input wire FM_ME_BT_DONE,
    output wire FM_PFR_DSW_PWROK_N,
    input wire FM_PFR_FORCE_RECOVERY_N,
    output wire FM_PFR_ON_R,
    input wire FM_PFR_POSTCODE_SEL_N,
    output wire FM_PFR_RNDGEN_AUX,
    output wire FM_PFR_SLP_SUS_EN_R_N,
    input wire FM_PFR_TM1_HOLD_N,
    output wire FM_SPI_PFR_BMC_BT_MASTER_SEL_R,
    output wire FM_SPI_PFR_PCH_MASTER_SEL_R,
    input wire FP_ID_LED_N,
    output wire FP_ID_LED_PFR_N,
    input wire FP_LED_STATUS_AMBER_N,
    output wire FP_LED_STATUS_AMBER_PFR_N,
    input wire FP_LED_STATUS_GREEN_N,
    output wire FP_LED_STATUS_GREEN_PFR_N,
    output wire LED_CONTROL_0,
    output wire LED_CONTROL_1,
    output wire LED_CONTROL_2,
    output wire LED_CONTROL_3,
    output wire LED_CONTROL_4,
    output wire LED_CONTROL_5,
    output wire LED_CONTROL_6,
    output wire LED_CONTROL_7,
    output wire RST_PFR_EXTRST_R_N,
    output wire RST_PFR_OVR_RTC_R,
    output wire RST_PFR_OVR_SRTC_R,
    input wire RST_PLTRST_PLD_N,
    output wire RST_SPI_PFR_BMC_BOOT_N,
    output wire RST_SPI_PFR_PCH_N,
    inout wire SMB_BMC_HSBP_STBY_LVC3_SCL,
    inout wire SMB_BMC_HSBP_STBY_LVC3_SDA,
    inout wire SMB_PCH_PMBUS2_STBY_LVC3_SCL,
    inout wire SMB_PCH_PMBUS2_STBY_LVC3_SDA,
    inout wire SMB_PCIE_STBY_LVC3_B_SCL,
    inout wire SMB_PCIE_STBY_LVC3_B_SDA,
    inout wire SMB_PFR_HSBP_STBY_LVC3_SCL,
    inout wire SMB_PFR_HSBP_STBY_LVC3_SDA,
    inout wire SMB_PFR_PMB1_STBY_LVC3_SCL,
    inout wire SMB_PFR_PMB1_STBY_LVC3_SDA,
    inout wire SMB_PFR_PMBUS2_STBY_LVC3_R_SCL,
    inout wire SMB_PFR_PMBUS2_STBY_LVC3_R_SDA,
    output wire SMB_PFR_RFID_STBY_LVC3_SCL,
    inout wire SMB_PFR_RFID_STBY_LVC3_SDA,
    inout wire SMB_PMBUS_SML1_STBY_LVC3_SCL,
    inout wire SMB_PMBUS_SML1_STBY_LVC3_SDA,
    input wire SMB_S3M_CPU0_SCL_LVC1,
    inout wire SMB_S3M_CPU0_SDA_LVC1,
    input wire SPI_BMC_BOOT_CS_N,
    input wire SPI_BMC_BT_MUXED_MON_CLK,
    inout wire SPI_BMC_BT_MUXED_MON_IO2,
    inout wire SPI_BMC_BT_MUXED_MON_IO3,
    inout wire SPI_BMC_BT_MUXED_MON_MISO,
    inout wire SPI_BMC_BT_MUXED_MON_MOSI,
    input wire SPI_PCH_CS1_N,
    inout wire SPI_PCH_MUXED_MON_CLK,
    inout wire SPI_PCH_MUXED_MON_IO0,
    inout wire SPI_PCH_MUXED_MON_IO1,
    inout wire SPI_PCH_MUXED_MON_IO2,
    inout wire SPI_PCH_MUXED_MON_IO3,
    input wire SPI_PCH_PFR_CS0_N,
    input wire SPI_PCH_TPM_CS_N,
    inout wire SPI_PFR_BMC_BOOT_R_IO2,
    inout wire SPI_PFR_BMC_BOOT_R_IO3,
    output wire SPI_PFR_BMC_BT_SECURE_CS_R_N,
    inout wire SPI_PFR_BMC_FLASH1_BT_CLK,
    inout wire SPI_PFR_BMC_FLASH1_BT_MISO,
    inout wire SPI_PFR_BMC_FLASH1_BT_MOSI,
    inout wire SPI_PFR_PCH_R_CLK,
    inout wire SPI_PFR_PCH_R_IO0,
    inout wire SPI_PFR_PCH_R_IO1,
    inout wire SPI_PFR_PCH_R_IO2,
    inout wire SPI_PFR_PCH_R_IO3,
    output wire SPI_PFR_PCH_SECURE_CS0_R_N,
    output wire SPI_PFR_PCH_SECURE_CS1_N,
    output wire SPI_PFR_TPM_CS_R2_N,
    output wire RST_RSMRST_PLD_R_N,
    output wire RST_SRST_BMC_PLD_R_N,
    output wire FM_POSTLED_SEL,
    output wire FM_POST_7SEG1_SEL_N,
    output wire FM_POST_7SEG2_SEL_N

    );
    
endmodule
    